PK   � ~X
0�0�  ��     cirkitFile.json��o��������V�wR�ֻk�z��p��,J�.F;��}y��?�l'z��d�v����6g��9C��ϋƾw��r۸���٭�����ŝm���,��m�����w��������r{��ݸM{�J2�%����ʌ�tVp�H�sc%�%���w�W�S�:��s����K����sʶ%��e���+s��F���\*^(�W��s@�R���l`]�a����q�@�)x
$�*����@��?�m��1 ��ǀ�1 ��ǁ�q ��������R��Z�9�ՠ������@�>o��	��&(��(��խ@uC�z�:#�� �3�� �Ƚr/���3ȟ��@�$�?	�O��@��?�O�S@��?�� ��) 
ȟ��i ȟ��i ȟ�� ȟ�g�� &Ο)SR����{}�_�\�*�[�JK�nO�ծs�sN�0�b�R���e3���-�U$�\m�+k��X��T3�I��D�����9vωC�9V�(���g��ꅲ����$+�����9�f��� Z�rJ<���pJ�H 5Ƕ�'O@��;I=�n'�Ǘ�:�l�n� X�	)6/�n�B������A�7M-4���n�B�=㩛��u'����y������Ǽ�r��6����H�X�(��b��X(V$���nVt�R2S�5��A���:$xq�8�R~)��`�p�h38S��iơ��P�p(f83���b�C1ǡ��P̑\	�yGq]�\;��#�ԇ�3w�V�, f�몐38s�Ţ�XY�T	1s��:7�#ƙ��\,p�b�3���b�3K��X�P,�;�%��b�C�ġX�P�p(V8+��
i�b�C�¡X�P�q(�8k�5��b�C�ơX�P�q(�8���b�C����<KqjΈ���`�V'	�������B	�3;(/Ç��	�Rs,����(5�!���}�
�c8*��Wp�T 5G�</�����M=�?���#Xyv�M>��0��D���ݬ����Y���w������f%g�߱I=�>�h��2?N3O'ƻֶzb�q���k��1�
C��Q�+ŊB��Q�+9uH���Kq�8�R�)�a��0Ł��P�p(fHs0��b�C1á��P�p(f83�9��b��J�P�q(�8s�9��b�C���X�P,p(H1��b�C���X�P,p(�8K�%��b���P,q(�8K�%�
�b�C�¡X�P�p(VH�8+��
�b�C�ơX�P�q(�8k�5�6��b�C�����Plp(68�ͳ'�í<;N�'�p+϶%��n�-��|b��,��'�p+�N��'�p+�N��'��!��C����'�fp ~��#������c���pY�_?��O߮���+ʗ����nֶt��js�m*�,��!_#�]�-!_�Y"5'�����[լ@5Cz;zωXCV^H͐�汚SO@6�nP
�li �I
�Q�S@�<�nH���*�O	$KR3�3�z���i-m����_L�[W�}����.Tj p�=ۀ���~��c���/��= \��6�k8 � ����:� B�^B��B�>�	`W�	P��l��� o ��m��j������>~�#d|�W4�����g@}�@}	�Dd���=1G#crv7��r(]`<�|R(�J(�"J��v�� j 
"��Ƞ$2�L	%�AIdP�D%�AIdP�D%�CI��EJb�A=Z6#�z*��^ĕOϩ�3{�u�D>]��e (�Jq�S=ru@��Ħ�"�Tz�5�����ζ:�
�l+��
(�ʩ�ζ:�J(�$AI�P%�D	%QBITP�D%QAITP8^����$*(�
J�����$j(�J�����$j(�J�����$(�J���h�$(����9ƣ�$�阜l<2��O�:���	���#k�SpTs3���NNc"9j�ɛ�ɹʣ���<��D�K�^�����d����?3U�'-����yˣ� ��:����!��4��A���N�m�$'9�M���#s"�=?�YU����߅Ԕ�2��) n3<�az�ahg@'w�Э�]�t��4� M�8�4(Р���l4X�`A�4X�`A�4xל���t�]>D����F�u�"ht)�!��� h��!��"h��!��2hȠ!��2hȠ!��*h�����
*h�����
*h�����:h蠡����ڠ���&h��a��	&h��Em)~��`z���������L��H����Ƶ��ÛGO��������zY*(qҘ��
�J*������7iL�}�_%a�J���Y�@IF��-�����{a&,p�|�&,7pҜ�ZMX��946���LA؋?a�����f������wk[�uX�G<������ʨ��贈�ش����H�ĴH��H�ԴH�����̴(?�"z�:����������~���m�8[[ۄ^����j���x�� �~����>w��6�״+����O��W�k���7ߠ������]��_��/��~��,�o��퇟6�{���ڮw��\��j�*���Z���_5�Z\��������}m�v߸�\�b��rHZ�tx�[����kC̥�K��K9��wgh����E^+�TƜ�Y.���ڬt���EA�W"?v����u��r�ô�nʃ��`m��6+o����?۫�\��^���%����Z��;�]��w]�������a��œ����w�<]���������u��]�dz�EI��(a��/���ps�ia�"�%����|�iZ:[��:*�#�:<�Cb%�ј-�Q�Qա1�e�%��J�������И��c:�DuTTGFuxL�{�y�.9���YN�눼����ƓZ�h�5�d��$kT�Y�i�D�5�f�&Y˓��$[*��<}���o|�D�于ȫ��<}�y�&b��M����E蛈��7��o"6O�Dl����<}c�y��R����KM���*xzR�e�]W�Y~�����b�oזw7���bUuW�Bp#�3U[�3��"3�2a	U�r�4��w�[�N���_�9�ҜW��a���]e�"$#�V�u�r�t������+!�0��3�&�\ٌ2^a"5�Q���a���Ii���L)����,�ʤ09��R^����l~v�ď�OnN��ӝ|�ZW=ˊP�������2�2�	�*+c�+��M�mzp�~�����*��м��󝑑�
'	�U�g�|���\�5e�T���J)k�Ty����)rZ;�����}����T.���_;~X����?Ŧ�x�xe�7W�v_�'L�%o�M���j�nw,���K��^��]�^�O���Վ�{ N�n%Ef��*\�jS�5>F�Q�2��a��2��*o�v\��T��V
���<+�C�£]x���($a�PY�Q-8+�TJ㫢�����	S��V���<a��ϛ���عv���?]|���\\������O�}s(��w�qˋv{��7[�\yi�ߗ�?���v;o�ޮ63f��l�����C�qkW�3]��,�rq�>�6)�N�;>��B@��U�K��V��xmA/�e������o4W�n����ͦ�#�4��SR
%��g�Q�ߔ�_����9���p�LU�,7�ӥ���꒓")�N:,�kW��p��Q���M��(f�Jƌ�$�_�󣸜�^hxe���!��/���}���] K:\M,������m#�C�Q�.sbdN�#~3��;U?����}�5Y?���m�m�i��R
�ss�h��:����G�r�GIW��J�Lj���{'F�U��8��
_�I(%�'l�e~�:���ܥ��/��O`jF����K��r�.�a��&2�}\�/cy~���_?��nN����R�\���|^,�Nx.r���-.�f��D���~:�"#������&��{��2򧡻��R��:5X�����vg��e����.����0�������c��[�:���g��M�ĺȸ�����V̋��1CN�9+v�|���Ys�h�P���z^n�f�r���Fsz�s���yO�Z�C�i��tm�L+��[K}tR�p���.����0)%�1�݆-7a[#�{�|7����~
'9�����v�g�Eƌ���.��[H�5A���[}XU�]0�9����[�v�v���+ٝ�|�~�e��s�w��Io׶�~]��
_�?���G6]Dp|�l��>mڷ��1�x���!z�TgM�e�t���̦y{�k��v�i�����僡�E8���~
~���]�zu����ۧ	<������*Ul�a�w_|��I���Ę�N��":At�1��7��1U,u��;N�����AO�2K�4-a�_к�0 ���Gs$��)ɾԓ/����{�1�<mrO��C�����{���C>�zr�ɹ!�HE���-̘S;K�lK䩝��Z�ҩ}t�>EH��w,����C�3U���Xd��^��C���h�����102�E|�?jK�/�"-5�[a����X���>�����Os�:�5B�i�Hb~9v`�����}/c��t��K3 c(���T��3A�T�g��ȍM��iS!�{u��!�=��K�F٫|��>d����0�'JY�T&g��|�T"e9�HY�R&)�^����U��p;��Hj��,I*��a���R���LW�D�L"r��9����Wq68�r6��F9K����z�^!��YHJS%*gi�:�����,yc�%�{!g���fC!��(K�������D�R����:�@!Rư)S���W�f����;:���g@1�Ҥ";��G2^*��Y�L�ט�!:g�k&�k��s���
q=ˎ·�MiR��pr�Z����kVv�[\Rv���sՏv�����oZw���}Y|�PK   � ~XWC��)�  � /   images/093f54e3-331f-4155-80d0-fca9fbcaa25c.png��	8���?>ҡ�)�T�9�TBC�,5��A�(Kd��/�q��2r�fP1ɞ�0�Q�
���=�k�}��~�z���������{����y��{�_���ǣkښ<?���\�����.��~r��>9��"�؉���]���u���K7�0ؑw�v7����0�='k��-�;0��v��h�[�wN;��ď�?��
����O�h�O� ݯ{~bz9a�.n���(��@�n�OoF�������_��v,ȋp�qW,��!��U�Է��N_�W��+��ޫ�}���.}�s�����}2lTSr��i�� C�s���sJJ��i%������鮋��?�������� T�źȜǾ�'w��A�t�+��OhEz8Ϥ�/e�>���e�%���%O��'�3W�L�����TV^&�o^����{��b0���.+Ű	�~�8�O�m���z�K��n��矌�t��d�D��`���JJJ�a��8�]\o7��N���;�Y��Kxrt�
Q����G��jm$M�KBS�='{�VVX+���i6=�˯�hT��_�1g���a��p�ݥ���6zC�*��4?,V����U�\p�{�3xc�w
C���\�"��	Z6�{��O$�O�(����Wj%�X����K���}�u�=���'�5�^%U_��~��!a�@G����1���̦a�w��W���4�8�$,䄞/���v�G�����^�-^CY�	�S�	�n���!T�17�!~,){$'L#Y'I�c�*1��9H	���|$��~��P�M�P�?%ͬLZ����{�OY�'L�oUۿH�H��������e%���OƯ���CkBW���Ou����Ƥ�n=`���C�\������Ŕ����ORŖ� ���۟��(����򣂒WP0;��e�*m>���G]�
�i�jl喨4eX���[\Hk��������6��ņ�\�B�m;�=��U�C�89ݻW���sv�~7%�f�J������n�2�oQ����u���^ۗ��% �5��£9�Z��;��� �1����p�`�g��7�Zt��nf��J/���DvE�.�5�b�`=ۥ��"֛�����K��ͫ��C��zCq'�sN�z�N�����j&ӟ�Fs�/��!�;�p�ԓ��8�L�aOǆ�{�����BT�}��dPTbߘ{1�K� ]���`��8�6JqSV�K�O���0�`u'��oB-¼�E��a��+��G���s�.��/�2��|cB��6]�`�2{��TW��wAR>ڦ�ªIϕ�s��}�z+/��Ra@�;�b�.NӍ�;n�`y�O�X���V-M����������D8`y��<�D�Z�5����`ҵ[���X8>�Q�+�Y�m�L�Cp5~"�i!����a�
���	�MO�����B�"��2�T7����\A�I�o�}8�àq�`_�K��w�.N��<�_��r+���>�m�0!��	�?���c]dkjd�9�f};OA���HGX��[[�klHR���B�I��N�-%=]�$X�v"ɑ4n�<���v�{Ы����1�����m��(�_?�'t_'s��n7�Z$qR-g�}�����
�3�U�	�ۉ�Bk��c�4Ƕa��?��d'L�_�� L'@\���P�>���u�y�f�O��1;arQ�	$|I�KՎ��^nKɳ�4X�,D�|��"93��"���$�7Y��y�������@�N�K�d�ct���}u-�D��g�w35_��e� �2ty���dM��E�Uಷ�'�;6>���X/�I��>�ѱ�*&��7_�~7$c[F�O-n"Y�'������N������-��C�*6g�uv�����'z
	��r�/@B����p�\j>l{� X��P���z8�&7/o_qq1��w�7~Gg� �5��O�|��Ijs$����md��41��=�Y���E"��ll�]��wӵ��x�aΗ�����b���w�{q��lO��5ޣL��3ZVZ*���L��6C2�\0��`�}�^,��J�t��B)��x�K��x������$zU׏׌<`ۋ��s�.���]�J��ˁ���#�9�!@'��q6���$�����/%e ��EM���ˤ�(r�1��zI"���� zZ�	�����߾=JM�>����WW�e��Y���9m[9L�(�������[��K���G---����f9�1{RYQ��&c�.E}9�]�Q���{K�r0?��%2�%�:^3�YO����?��dH�UND�k�@ �lz����S�9��Fp4�����h�]�|/�5�_DJT��'A�����^AW�H������ b^��z�����z��efeU��Z�D"��e�wI�o���Һ����%!��k�K��n�^������rs;k����W�+���Ȉʷ��o���MI���Z�]��󘻕���w�C������FF�@s�F�j��[�,�HZO+�qm�n���@_�w�{����f���w�_��6r^�@�I>pC*�ӱ���q;۞=�)�@e�A1�E#I���+k^.uK���'jM?f9� 8�� S�@�T��.��w�=��U]dnI�p���{��%���kS_���S'(,�Q	f��.�����f�kn|���Q�+#��
 ����g�T/�����Y�y:a�x�[�%���*����f�4UQ@!/�2��p����W'Xk����u��ӧ��e���[��S��7��c}:[w��1��rv6�b𾿫�a�g O^k8��<���f�\^c\�s0���Uv��w�
ܲp��V^w�� ��;��?ݨ���MC� �M:�M� C��},\K��RZ�B�&� xVZPp���X�{��E͎�Ύ���S~�=�y�tWj@�XV ���<G ���ؓ1�;Zv���5���Ά�V��l��&Z�	Jh�^��kd����o������������{珰���6�)���i�,w�&o�@�X$Pڡ�� �4���Fe�)<�8��O�!*7141	u/6U\�� +܉i.��0��O� ƺ�:w���f?^7�^,sp�f��t��lhf������8U /���@����l�T�	�5��it$�ޘ��%�O)>������Y{�h���t�����	�m�ja)P<͇]����(wY�o-yꔧ�Z���x�[�'���<��G(�mm��	��X�����Rp�[`)}�ROG�H��F�E�8�3�	]��}��m�L�Z��k}�ES]�w�hA�r�����C��ќ����.�&��-uC����|7˴{a֨��fvXq����Ps���<{�#S�Z@�S�d2����U�%V��ә������q��������^}Avֻ�s��j��A� ���f��U�(V_�N��j���3E:�SO(7�|0��5w���P\ؿ.,<�<g���� ��Fe)�X+H$���4����F_YLb2���D1�_ל��.
u�ԩH���gv/V�O*����w���AS'��EA����K�W�"i�Ts��_Zzz �XPP�'f�V�u���7��:EvQ��~��}]i�Z���{��oG�+��C�3�p��HF?v����;<=�Ez�����&[���j�����$]�A~~<N���ie."��Je���]m�=ɧ<���B��p[��k(���Z�g�_ou��Cj��Z�7�]��:�/EEhV�Y-6��L �W�u_�X��M���y��J��z�k��/-d�!B��������ۤ�3�6hBU��]��4�,��� ��%���^�B	���������6�F���ă{��lp�őhF��Øq��~�,�G	�k9-WvĢ��p�@SμL]��.�bU�T�99b���}8�u�HrDq����\��j*bcku�M#�� V��Rh ��qprR�z�"��ž�AQ��ĵj8�}}�EW�#���}l�<&�8�Q���xr�wR��`��Mӫ�
�A�M��(ƭ���M���o�������)+۞$�ƶ��J�%%E�]}SR�;j���oԦQx�])== &8�����)�J���u�rY�o	���Wy{��_�r ��Y��=�6�WC��U��<�f�i"% �k��3r�"�zC�����gC!�,�J��b�~�����������n�	�6tBHB}��z�����d;����8GRdg�w�c@��
��l�����0YeNl{JJJtqեӭ��d����(�ȧ�����tl�3�l��vd�gS��J��I3����?ͱ���6m�c
^S��IV=T���ODy��t_s�V
	�]���+�}!h͟;Iv�f�B]Gը} i���4">�)tf����<4��:��J�'e��-�([.��z��.r�)��M�o �0d����wHGܚ�/f��?�T������K���k�=�����o ���>D������C�5a�]���+y��_�������9�f��*�;ǃqX�U�^MO�p��L_�6�p��͆7S��> H���j�8}�N� �V�5���ւZ'��QH�������9����Lv{�M5���;�]:m��{X�yx6�
�U���ꦭD�X��l �@�T�D�)�]��<*la�PWo���ux�j��rF��!�Ne^p����O�̸�t����_�YC	R4���&���JJx�Y�.E�ɣ��S���p�j�T4�J���қ����g��.�Q�'���E�'�Ν;WF�삭Q�f�j���1�6���ک�<�éQ� �e$��ݟ	Z�Ys3��@%�-bz:T�)^�/��~q��SfK%�/��^6�ʯ�$�DY��� �O�5쳳�SF^Wm�+$Q��\n�$ �k��#؞������,��I�#����@+p�J�Ȭ�>����"̎'�~�����o�ċ����GX;]�z�@�~���&_֟˝F�49��Tzϒ�V�����Y��s�3�g��`,�H���k��yl�=���9>�745M����j��Ry��w�TB�M��	~�[� ;��`�h<Zg��~�v/wu�4����6Sz���J�$�ZҕђH]�t	�訥#P�>]�?K�����V�Q�;-���RampX�Ř_ާ<Q�hߤr���R��t�lΣ��D�Pܪ�=劲�|�������e�]��cl��֯�R`�,}�6]���.��Wf��\+x�+��W���s�Sk��q,���Xwi�Fc���}Y���l(��+��O$.i2P9ި��҉0r���#�h���ȁ��co�M�͡O�0)�J�[��� �������𝮟���S0x��1�a�tB9Ɛ�`�G B�KT��Z�� ����d�|I�u��]jDؿ���*@���v;�i�U�2<T�}�rjk�e��i��������Q�+Aw�&�e��=|2;�����R\Z]�:�$��@�%�1�z۸YV�(P����Ŋ��],�|M�G"*��q�j��r�J��,y�k��䐐?�#������������&Y�]^U���3�8^DO,y�w��\����>V�<߱���(�@�ƠQI�k�,�س,//����,?%��1��˫h�g����Է�S�Q:b���n�s�{�wͼ\h|�"���I��)�i��+D츷��� w�Ә�i���kÈu��u`�����$���v���-T��T,��UE�K�X�Q���g�P�A�fؙw��a2@_��5��8�'�fyՅ� �"����ay]>�H��'���$��[��
&�Z��}��*!Hu!�s�x�h(��ݾ��. h�P�s�*?��_�u��Nm�ݝ�~�C�V����������W5S���7�x�L��h��TE�|�A�����A�#���'��ݓ4[6�Uno�vB09;���L����;��q����d�I�H^�77��7o�G�z����O~Lf]g��&+�k%}pM|$��KM�'c�Ck��Z)G��B��Nii�E��ih~X��|�~v�l�r�M�����J�p�sM����bta��I*���f�����\W��,�c+$M���g���Lk���6;Zq��ɓ�c��m'&&X��o��[�VL.��dc�)-���%���w<���n:���R��l��H�cW��)�M=5��KA8�{��Lj��r���s���$�}a�֜_�  �S�O��w��>�ɂ��B��������5R�Ua0B��[�2���Qq�9�#�o߾eZBlL��o����/ �����������X����gO�?�7���_6����j����H	�xr�M¹�-g����3�ƿ1(ZӨ��i�#�X��IYQi��(�@+h�X~����pG��E��֚�(TU[�ԂH�}���S�F^��<?k�PEU"=[+~�C#,�\����RqQ�M�\�O�0�
){Z�5_������֞���V�i��mvv��	��bd^��I�ø{n�x�|��333:P�����A�p����x(ӎ�����AqmN;UO��	j?p���|`�g����� 5aW����'?p��%o�
MB��ϣ}�`FisؾȚ�7����nM�brA�
�	���/t�2¼}��Y�0a}$cIS�o��t��R�A�(�6���:��� �<J;�d�X�bB�xZ�ܜ�_�OhP���=�oI$-�p1���-��'� �"�(�U�	]����^��9hbs����ؐԶb��:%�ؖ܅?���A�TS"�n�i�'
�P76+=�-GRr��fjs�U$�~0�&��X ��KӻZ�>h �q@�=������J�λ:�A	����
b�<� ���ݹ�_[|�E�jf�)I>��� ���U�h	$?qq������\$�[�W�3!�d�&<f����Ļ!������~qm ��6|���TLX)���<��Ьw�?�-�x� �1 ��!_���C�p�r�~�M})�y8�7� ���;;;i7����h���(TPAHK?��꿇+�U:�|R�(��
>8?]'˞Kwu�12�~��Bo�m�C�O`i�;��@��:نJ�V���#1�!����>��2wfD��t���^��s���0"�Wh���[�m��W���-��!�`��gc����ŝB! ��84s�*��IQ��@��8Ȝ�995iz�� ج��\ޒ1��o``u���o�><���[�hȽ�����M�v�@Un+|��Ǟe��� l5�ѱ1���k���aY��T78VFy�����/n��R"�k߹s�#Z4�4�R���c[^t�BF�wS|�#I�n��Ѻ�)
u���T'S�6����w�0� �����/��h�>nAd������?mP�}���M���㝅�@F��&���{{���e	���Yb�����A96�	��='kYq߶נ�2��7��(|]�_��J5	�Om�����r�;G�����fF�6�]��+֘��}�H`����у������O��(t�?���̗���vh�
��2��/��
Ƚ���p�߫�NG਴CU ���{"��`������z��7\&;{(�t�u��V���D��+�n��SRI��R����n��}��V�翐�����2gA���r_:p��(� h���A�@�5T��.�4Y�St_��k�ׯ�����`	���F�s=S�a@_���ͧl�����9�k�f
�{2��Z)pڄ�"�<�ޅ>����% A�
��i�t��rmSu���QI8c0TT���w�}g�w�燼*�
��]MG�A�(�q�F��IԂv�<'��y�%l5���l���b�V_�P'�K&��!r�^��%�}�i�}�=%2���Ջ]{_dgqx�>/���TF��=���+��z��h�s�n���w
��B���u�:dt�P��x:����ms9�k!�t��Y��n���c�p��ۭ���T�is�-���R���w�@mԶ=�_V\�x#�[�-����������`�ݸg����@�b˵- a���}1v�bon[�]��_���&, �b�a�7�I �Љ��	� ����
����䓟�1j A7Q�Y���F���Q�(рN����goG//L�a��� �,�g���:8�uX��7����{9x[�?<�z�>�/~�s<�?��m���Y]�5�/L��<�ǲ��o��oT���u��������޶G�8K�6�.�f�l�W���t��Z�~���~�F�����ȝj!�FQVgdo�S�(��(���y����e�D}z�CдI��Kg�˶�I��k���/�������ہ���@���o��ÓǠ�`y���
����}y-nVm[qLbM�����A&)�9����I�������.4�՝��WĦD�BzDm���5�֗�.�k�����z�e�� Ɲ튌)(2����5�#=@���S���hZ0C�O2VO#�n���K;�T����\�r�޼��w�rq���Ѭ��e�D[�+�ڶ����qO"M�-<�}���L���]��ҷٗ�SH��^��ČG�2�	�+[��H���7���2��;���S�mn���4�͛�O �a����.<���8�~�g����gB���	�׹�N������oR����,L����O��Z�4{��/�%on���3��E��Yږ������:�z� xݼc�Ti���%���JܰR g̚@"=�o0IB�b6l�켖A� �8�z�#L<ՈY�:ѹc�aa��@\˨�V�{m���n#V��x��>���<K��au�h����d�gu�;u����8߆y^�"��@�`���T�1;wI�/Ok���B�Dܐ�����_F�z�!M.��u��K���r�%��OV�Ն�*���	^��~�sbp��&Ӊ�i�B^Se�}�q ������[���81�ǘ�DM�"�D�w��Sp���G��D��D�����)��4�T�����::2z��� �1/yN��1i���3�1��!�!�?"񗈤��}8o�5����5(1H�(��f�����K�:���r�W%��TWDۋG�(��^g��º95�dro�N�Ж
�
��D����!_语z�X~�F�p"�^�h4;z"�&52I��������F#%[ \��Ng&uY�u	3��UR������j�Cʴ����kJ���5�Zn�W���O��T\w�B~s[��r��h�&l���U0�ъ���������u=����(�W����FVrp���o��M�f�-��{_�:/�K*	��	׺�l��&C灧�������}�����*���j*�uը��ΟF��1�_0li������O��2B���U�e�St|��_�m�+��;/�N���L�X0���U{�ét�V�Kx��,|��/Q���W������NiV���)��;�TV$&X�q_gʗ��Hʝ�~���{68/'�^��������RC~���p�LnE�����bt�%���qF*Ӎ��Z�EK'�7�\<-ֻ@��ef(vu��ZYmyB�'_���Ǵ�3C�n�S�O��J�H�g�B4����,�����n��ު҉���[� �=2�&�mU��}�����_%�)��	��U�;����3�qY��d�OUg*�?:o�\S��w*9�Zx~ �q3������%��r�if�W�x��*o���R��	!���)7�/�R����Z�vJ�az��a��V���H��A�\�~��Y��vإ!<ĳ_wΡN%f�W2�>�2����P8���`��o0�'a��_3f�P�h:W�6�	�(�k�2v@5�?�4��pd�!���X�����VB�̡���&U��Eդ�(2S�?�McPi�U�2����5;|���&�-�P�њ����+�����4E\������//	o�+�Ӕ7-xj ��_B�*��f�/�;�yd"y�S���Ā������1�q�ܚ<<��Z]ɧJNm��ޯG��9�1 �I��i���U����y+���Y�j�;����307MU����#�(юYK�����vO�h�x�S!񥘘��~��WGK����>
��$���m%�JB�҅x9��f�g�%�iz���8��-���b���fi�����u˯'Ȇ�/7=�ߤG��i��؊I���6��ϴ]jiӸ�s�_�ߌ�Q+��<3���8sO��ȧ�ZR�7\���q�c��*q���sZ�����G�_O!����5~�z�Q;)w8y��Hd��O�o� ��9�S��&�v�`^�� ���q���	�#�m淪��[�>�4ɼ�(�$PwA���� &�<H���rƌK���$� ��.zJ�C�G�m�߿/�3S&�o����^Xs�>�t�k#�}V/�\n5����X�蛺4��)���+�:�6���������¢':7����蝈W&������H��ԒK�E��R������ϻ�8��\W_�;Ж?�������;��[�B�ԩ�)�Z���R#_�g(��dgg����S·"�O�i��vE���o�����!1�1 ����k�_#����{)w��-!W^J� \�#��#�EEýK��i�=��/]���xxh������i����[`糼�^�o�0�LMIe��Q���G"��ej�I�:��j�$�]ۓ���QQ9~\�i���8,6q����GDD�p@�Ѯ�Vz���сJ�c't�U�ȫ�Ȋ���ݽ�|�U�ik�x�u��]XEj����&�ʡ!���P5���p��+R���ے��(�e�Z4�@c��.���D~e�q�#պ��N��>!���n-�șH��<:�C�rr��� Ä���_�E��'�L22��<�>>>Z�� �A�a�X~�b�S~J��z�~�E��L��-��&V{�Aȧ&����Ԅ�W�����.���_��4d���zx�ė�i�ɬE$�D�듹yմ��x�z"惤
�4 =dm'Iihjj�^��L"���T���nH���{%a�T`9�O�R��7Z^u=�U�+db��C
����A��6NJ��=����)4,,J;�}�[yn�۾���p��U%^�Hq��CPV������OR$��mR����o��`���JC��-�H�u�B+F��Ç6��ꁷ=x� �,u@�L������ᝃ%�vmc����c���O%8t���������^?�����کS��[>
y�F��25���hW�ҁ�&
�^��lfC@Ǐ���W��;�|H��ڝ1Q|V?ʳ�q����9^899���Q�U��}�����2��3���v�^~(����&���j���v��ỒWJ�l���)�cv��L�>���H(.X}$w8�������`"$�B��#w@(��k>�cZw-��"k�����bm�%h]�E��)����ۿ�ل+�У��ī��-4����5I�Y��tx�+^'ܔԜ�4S%4�5
����l���U-i| �L�����ӻ��[�|0�	���c����\v���ml������3N�_��Tg�H�UY=����4E*��������i{.^FZzom�dHYY켃k�<��v*�~F8m�W�9�4���1��o%9AϿ/��z�Ds8g��,<���z���4�A*�v�!P��}A�!2�Ǥ�`)s>�7�����W/N�ʥ�:��`�5Oԇ��ntGC������^����T�������C�����R/�@�o&��k�B��7
��D�7��[�tᲄ�)䬧�|�����7^5���Q��L�ʕ+�==��TL>0Og��+5�6B����̺���3��.M�ូk��ϯe	?��9O�o�f�7��j�MҎI��sc!��ă�+���/�<9�~�5�+y�ٝO��3�[;ᮊ٘�j6��~�o����W-ws-��E� v?�[e�|���B~:�~8,��*mM2���j��Cg�(\��H?i�C�v\�+
�#���xEnX /@���-����W]Ԧ������ˊg4����?đ]��=�{+7:��z/�Fr��3�>��@m�����ſ��E�eu�9^4��l���V'��s,[i@ἆ��@������"�B��?<||��fR	2��+[���Ow �pRj��w0_�m+�vu�-+�i�2W������ye�z��g��Ď�I��KO~���a��WJ�yp��Ԩo�Y1��`��%2��Ǿߴs�=�>(�"�	���o��ci ށ;!m�.�J��e1�oAߪh��0������a)�.�}���I|`�(X��8��EO���&�0zéVׄs����gϞ�
>Ua>�g���;���VU�����M��BӃ�!D���7wj-�����9�K[Թ;�U^�	+� _�q�X�AX���\Y�mydW���o<ԏ�>�}�z�jk����-�!�6
5$�ғ�T�1�8����"��pE��Ґ�`��eW�W����ŋ]*�5Ր��iqB�T�2��=���f��iiJ���z����&#���/���[��t�8��M��h���#4����Bv1�py�85�����j�Qe�ѹ���t��FE6q��^%S#����56==���S!��M]ş�Պ)ȝ0�k�B�Wͥi��2�u�`J�篢���w�J0S0�Ƙ8]�gnT"a2vy���>�q�{u��f� 0�|Z�ݠ�k���0�R]أå����������N�i�c] �02�	o�./���q�i���ʒa��4悙J
�Sh{�b�l�Tr�5�����dIř�W]�����bk�@i��4_͵��+|�{_�bֿ�ߑ� ��jqj��[Q�K+s��AE�M,�E���Gj#\<����0���dM��ORV�bJndE[U�����<z�h�A�/@&�~B�[Va�X�>�n�mE	�����:w� ����d����:.��C�K�:t���K0�����3k*I������Q$��󱀹<���V���R٥sm_)Xl<���QU��^Ԏ�� R^�,g�[���9���,�J�YU#�b���I�dA�;k؜UDh���F����<3�<��6�;�G���n��$`F11�**��d9�%랼#��X4���f�;��86��4�IE�A�to�����k��"�4�	�E#X&S �T��鈂�j�����j��h���¹6����� ��	�B�.O�-�DpܕY淼�/�����߅�' o���h!�A�|������O����m�h����v���1�l�I�72�m�ւr��� ���A�4q�vg���/e��?@�k,�ȵӻ�����A���3Q�w�Ų��	A����3�{yL�5zE�������rT�����/Y�}>��fZ	����\bW��6ߦ��ʷݎ&˙({Ǒ�H)�>�'@|6����a��E���Ϲ�X|�AW�m`n[���;��Ż̶��|��S�Ar;�Sr�
coǼo����щ��]X����og)ͦ-�8a��O
҈ޫ��g�����|eN�K��%��ǽsg��P3uB�����V'H3uqg��&.� S������P�b��%�M(�P�#R:��m�"��j�I�<WU���d�WWpŃ�-���ϗ��r�\ANU�Gw'M֦����}�c�O w1+A�m{��ܨ�dNz��D��D;j�|�?�����$/:��4�d���������QN�ϴ���Dp�FJL̆mJ��׃~�����5�ة�RN���
����A��j�F���A�e�epϘ5�H{!����]�����"�&z!��#�1�/��ѲL����k}�F����KJ��'�K�c.,�\ ��'X��>@|�Jy-P����q��BG?���(\�j+o)��,�㥩G�LL���qI���1���t�9B�%�Js55c���V�<K�R��H�"o��E��B��zsZG �7r=P��~Y5d�eU�Ĩ���G!�i��P�J9;�7-^.	K�Vݲ���g���[=A+v����|ױ�A�7�o
K<iw����:'''@����4+%����U�h�
�n�T�?O:)��U�-�}XT�Ջ���4i�_�}�k�$M���2J���i~�KX��Ț��$Kޯ�$�H��t��+[�"��O���r�xaԾ�����M� �h�H�'�,KF}�Ň�|��kj��+F�í\oV��+���g��8��(W[9.w�^�5�Dݝ|�ar�y�}M���Fg�E��C��ے�S��.�����ch٬dNNN~@h"{�ы�؃!���e%��_++}��$`���i�J&��t���.�4���_X����vZNR�>y1�iL�!T$^w�'��S���\	u��ŉ�!ϘZtG�4b����Ȉ9�;Ӥ���Ғ�J�w� ed�y���a��9=zd2���ZZ�6KԠ�H�{#�I���T?98.)D�����J�s��sj�����{��.Ȋ�W*�.w,����/���A����B���͜Mjƃx�*M�F�4�.���냺vtl�@�'IY�B��
fw�u�neC�X�:V��wv1���쵻������G9��W=A�M��q��-F�N4��������Y�ң��VSID�)@v��}�+x��F�}��=Jfe�1�.�3��,�^�tu��#��w~R`�W�WAAA����Š�ڬ�� �R�vQ�]	T����6K�Ɉ�-T�$/��<�]�Z�ዬn��IY�?2�����!B��e����<��RDc}��0�)���볁	����>͔H�z����݈׋u������n�(T:q��C4�uh�:�CʩM�u���\��.����g��"��U�!(�����Vۣ��0u�L��Or��Ԡ����~(��E�]��>?�i_��r�k�w_����(F�.6�t����'��(k�X|�o��꣹��A/d1��b��qMh�԰�ǡ�
�\��#N_�?չCR� �E~s�2U��"wl���E�+�_��Nl{�����s(��<:���2W��l����<�rW)�8���D+V��*����Y�� ����v;!1:�0a}�؀�X�|��U{��n��k�j��XYN�p�oO�.��EZ����]�B�ռ���uv��&�3d�5��+�����\��{��*�WEn?V���d��k�8x/U��@r���>Wo��@�ӊ=!"�ǫ���o�"/��(ned���7.766�&5]6�d~X����Y�ߗ/���m���c"9o��d��"�1(�A4�= 2� "E~m����ņ2��AYM�OX!�u����Hƹ��e�Ӈ��V�q��7�1�m��W�hD�+��B�=tas	����Z+��l\D>��-#�=o���*�0jݏ�W���_�]nr#��RQbce�c���Y ���\�:�eu�ۄ���?$ٹ��?��w�Q�0K^�L,&�e���%�n&�7�&����f|X|/��I�����1�sf�x�?�v�Ӈ�m	�e����~���@�/���$���Cm�6�G3��Q5Z�n��� c���������F��V)�Ŏ��Ģ�����9��bE"���k�j&�w��cO�K�1��W�'�N�}HSUw��I��|�%z"ᬱ���_:���u$U�Å;�(V�~�Nh;l�X��Ԑ��P�F�YxΉ���S��.~��*��	Ct�8�2��s�X.j��:�^��2E:aO���R����a�T��Lw'|�"�l�i���gɵ�x��'ѣ�6��FW͜qd�F�i��������x"2�5+Wh�u���Be����I�t����9�VkjMt'��V�`�(�@ݻ��#D�:�C	�4�
�:���=4�N$T�>;�;	O�����)0�>r�����+B�!�ETz�gS5����)/$P	��&��d�;.?�;�B�� �^�_˲anL��)R{�[,�+5��g�..
wSn}w5F����9�:���u�q�%��SV��Yw� �,b1P0���r%7�&�I��5F�uZ\W�����6u���3���4+�76��,�p��O�C�H�x�V��[�>0?sz�Ze8� S�l�jh�v�@"U�Xw�����S�Q����g{a=/�}���É��R���=Δ�/\�g>�`�s����Y �_���.���氂>L�ý�r|~O������d����Uo���]�+E`��E��@oյ��gJ�@��F��g��!�BWz��L��m:�6�~�I���
q�H�.]���y�ń��v���N�����y�� ���/L�0}`� qD%z��,�r|RG�\pĖ7���yN��L��˴J�T�ӝ���)�o^S_F�j6�����$�OƎ�B�~$��E����a2";��T˓�,�-��I�Gx�b���i��1U[�d@~*��Ŷ�wM��gU"�o
����T%�O���F$���	������y����'���e�|
^�߱@������k0/x#<�g�}�O;!����3���e�0r�I-"���/��Ί�3�>M�֌��>��r�,�;E���O�^� J��!�m�mï��Ὧi���䊹���W����RԽ�r���/�%��^�d���v���K4�w�n���Ga�wX��dH,Tt=u��O-_Uץ�����5v�l�.ߐ��X�u#{UF�Y��1t��'럯���:�T��ax6Y����!��Q~�`�	�1�٣>�m�Ŝ���j{;>�
Ψ(�;g�Q���t��D�^"n�2�V�}��1 ��Y��VU��a�yNJ��(ލ7��V���5`o�����_Ƚ��Ӻ Ü�rk�0f���Mp�ծ��U��2 ���jK�+?|HIo�21�G`� �5��}�Ŀ(J~1��I�m����V��j7g��rY�|2�M�s4E/����#�/���8&�4�h�|�xV	;0<�e��4t^H#����Ǥ�)zƫ�ٹ'Rˎ��o��!D�T�����_y��S��&^ܶ#д�%�꛻��7;^�`�V�z0Vy9^�6�uou�rj�]"�(�8�V�V؇�1��������}!�s2l$�,���ů�x���}%q%�zl���*�qg�>vr&�i��[��5���_|ഉ1��U��&��ZϠ��� :2U_?��� -���	N�{���ݯ>��?���'��~Ǫ��'���A����E+S�ޑ��#�+�)0{yJ�n��%z����8�����x@�p+��ƿ˹\����8p쎎6��^4�F'�w�cO9Į^�cr�%J����^�~��vz.{:��f��9�St�J
���#Le�G��H�6z=n1��o�`W��+o�g��"�<���F�[��;:?U�� �˒�|��SRxv�y�Ԭl\R�AJj���nN���(rPG`ަ4��p�ʤ0h0��px�6��§�`r�u�����mv�N=����O~�)r���e,����.a�����O�/���W����m�@��3K�W]-١»�$��ړ��$r�nm��B<��k���'f�إ&���jx`&�_�R	݅ ��٬`�p�C?��=T�=*��$��.Fk�"��#
tJso�?9�j�y~\��YX>mR�i(�ab�A��� �~�����C��9,\�t�)���>+bƺ�F0R��$���+q �����Ҡ�!
��6U��i���vI��Cv,L�RlU�EK���X�e�o_A�~�>6�ŏH �Ib(qTrI�ɶ�FX��IR�\�u�|�x�ͥɁj�1�-�a����h:��������,k��AP!TwUP�"]QP@Z��J��KG�zD� A:�C�	=@(�|��Ͻ�����������9s�甙9S҄�{�|e�A %v��=3'<�9U�ԒN|ќ�nM��XbہK�ڃ��,�ӑ
�w<7�6�׮�K�~��-��g�v�Ս]0fgVQ.��{U��yt.� � �w�v�h7u��R�9�?!�:M�=Q]k���ء��;��� �(�� LYP%k�|g=>J�ܳ�S�0�a��8>���p.��=�õ�#ůY����Z%6�F�Y#΂�Ne����<����u��S��L�nt����5�D}݂Șm��Ր��x�{a�r�ܿ�V�x�ᖅ/�v�J�]����h���bz{�Ҿ��E����
o/i��������H���k�;�}Иn�Z�oN�����8Y6��9u��=�W��c�ly�ӎ<ǀr���3~0:^{��Pm���g��=����Q^XF�.W�����~��ǈk�+�aG�8֒}hkMT��s�w_�MI��m�VaQ)z+x7�Oo��Pl��q�O��W��6�ї�)|V����a=�l�Pva
��L�-q�#��)�{R0\�@y�Yb�0x�u�E�/�i�#i�|�k�b��tJI%�RC�?w�^Xn8��|*������'�-�?�e�9<�fR$4�V����<������y �Q�%@�q�Y�'�k�d�W64[<����ɡM�eȺ|�r�E��V��W>%e���y�:yczcF4�����.j}������n�31}5�,�X�d#���
�!P���+o����ہt_:音=�]68E��ˌ()�������<Fw�^�8.o�5��:7ݙ������K���LuV�_@x�����{��M��aj��⮶��m�2_lG]�)
�(��	�ˆ�alR��#r8�:S��%)?:s Ko|�60�m�۟-��w$��b�#:K�M�MIzs���BӡBߵ���=p?�N��`����� ���8H��j������~$IX�n�\<[���}U)CX�'��e}4T�Ua$��@��I��mo�M?�W�Ś����Wjn6'������IԄ��FX���f2�vY��>z=-C�ֿ�hH�I���;���P�:� ���n��Y���ys���7cx���t�E?/H<	�P=_M$)bR�����HC_J#wZX���SPJ㨚�a�v�!\t�"C�ѩ`�t���3.S��+��!�}1ݻ�m������lA�g����O��*Y��Vj.��M�I���P��R�;�hv��a�f���qC@9[�3����?_�����)�O�B���2�-�b{��V:��P�g��a������� 	��"��7�F�ﵣ%���_��%-�</�s��X�әU����K �����8���A�J�Ջ%6j��T�R;�]���}�겂�<*��[��I��sk�U 2z��v�7G�q%H;��(	V��K:}zEtRoo��8y�;�Bi*�(I��g���w��/�]��~Bۖ�f�ҞD���G0=�&�[�.)u�"�.c� ^�����$�i��@j�M���)_KP0�gl\g���iEԶ���<��9q�w�R����'߶;��k�bt>T�y�|"Q��8�B��E]���9f�ze���4��V�)�#V�Ћa}b����(��.?|b����A�ɬ��ԑ�%r�
�(�lUGR/�E9��.ٚ��y��`LdfNE�`��>��RV�>�U�M�p��M�X<�j �Y�)���6���o�&�0#J��F�MS�eE��K����4.�g|"099y���%[I�RY1";u�'�}ݬOW��nʤ#��})6���,��V���>S�K.�k��Зn��􆧚q^��.sX�qFb��p��~L9R��3H����k|�m�<�N҇j�jSw�l��Y�:��-!�gn�����m��E��_hL�Q?Nv,�k�M�!���]��=JT�w�?~����~�Ѝ�dy��*_�����2��v��-t���Cw���V>��R�^�a(VD�4�Z��]H`@23�p=�v\I��
�._��JܸW���γ)�����i���b\cLL�P�m�����=9��X�
��E6v[me<)M@J�^��Q\�ѣ� ��~~���ZL��5�؂N�ϘN����-+<�b����l̢B�{�K�;)ʊ����|�ϗ�{{{ێr�!�h�u~t��1�.�9̖p�y�ISt�)y�Ҥ�ECc#2&��C�10��{�j�ڠ��_AW���rx�0~-PIF�L-ʊ���~ඨizL�J��O��߄y�e�~�|�ZDv��*�%�:n�Z=v�.�-Mb��!6=�ĥ��g�2��vٕ��v�����Z�U��T�E��^��gWl�{�J-�s�����"�Ss�,����ﰌ��mD��aiR{�����N�T���-$xת K��z�R�Я�_O�×	����XI��HF�y�=)Ob�
Q��UJy��<�*���G�N�K����Y����j7!�R����V��0�;v�x�R���T [�`���d.	���P�fj��]�c߭��?��,V���������,g�lҚ�(���˲
1�mé@)�'�:/tf��z��ݼ�������̃�qq+Þ���������(���j����{
R1s|m+��a� :�<f�Nuܮ����!�Df�"8���W���~'��a� 6�ˇ����~�+��B5�Y�u�nP��ľ���N���(����OjM�I�9G�@ny���&�`
)�j6N� bj���t�]|u�E�L~+M?�l�%'w�b�'@SRT̗� (�h����*���������;2 `����zj� * d�v�i11��:�u������'��6%%'�*�d��\X�Y)�S��V���~�\3���"���@0� ��mT�d)����;G��TTT�f{r�w(�>�<6���c�$�e-4�!��e�j�u����u�]�����Ri�-�����1---�E˿1��z!4�mj�>'��6� w�yH:|] B ��(����4��~'��;� %�u�
�	;�"�1򷳧�[�s
��iy{���B�ҕo�k-PY!O#��l �-H�2�ӵS�S@4q��an�KP%����2N� �̚��Ó!��7��Eށg]��3՜�Iq~υ�~ ��	X,�y�Ɨ���@����]v#�������_��� �}��J�j+z�}ez�ʂN�a/�$$�iX}�O�w����d�Ӣ�dM����r �Gc8��ٯ!��.�����_��	�Ċk<�Hŀ�7���5�%P��,�ɒ�~��nw�y,GQ�^f����ߎw1-mhԎ]�z��`@R*�Ĳ]�E�	8z�x�I�w��X�S���o�j�:�gg�n��o���
�6,�ˉ#�ހNr�~�E ����t�t�����U������\��"xSy���� ��q8������v7�����I�A
P�/��-���N�ϱƗ�rp�q ���#K� U�������m��{<d�o�h� ݪܴ�yW��~a�:d}> ��v��@p�5yZwY]��1�m44{�l��a���i�D
��ޞ����iu�҂���֌1�;��-d�
f��t��n�o�W��ٞ���)�)j��$��{ZZV����Q����Q�ee��s�v����ͽMH���אZ)0��s;�L�4��&�ᄄ7D��9�IK�����(Ah�7��HڏݎE8����}�^33775������	��V�����t�?���n��.J��`�1����� ��m(�ܞ������FUM(�{�!�x'KP�����k�#��~�T<��Ú6��F�d���~��	ĊW1*���Ħ���X(�.�HC)�E��c����\��8M��A5�w��FgO=��dTP��6m�2���/(n4]�����LI鴨	�U��&�]BA9��ʏ:^�A�O������/�Q�8b+�vnJ��K�2���������2�Sɡ��8�BP ��2�#0� /��h��j��>���SIzJe��՘fh����/���اW��z�"���N�+��?C�+�m��b�9 ED7�G�H\��(�6F��7�ܦ�����v�C�Pi��|�d s-��a�r�E�C�\��ֻO]�����/d���n<謥���*����K�$e����Z��%\���6AqǾq�G!t�!��yw�	�|�Wfd�S�<��9q+4�N���f�MFW�G�:�?�T�}k��u{�4�8'��� ����J�&
&�=ؕ`��9yy���S�n@A����G�Sz���8G�Yo�ԫf�h��@��h�kV=��_��UH�'��r�H��I�s<k�lKb�:��	��(V��CG��b� ������k5X��J9�?����JA� �*~@U��0.{�0{4�}�h2)Z+��t�ڻ�C��淎�yQ�2���p5p#��h�����ڞ�.�Az��
�#$��j�`ٮ�DC�+�޲�v9%�<�H��S���Cϡ��8-��Ժ�U2�nh���e��
+�P�9 �@�߃Hw ��{�@�����d�׾s gM��R @&� �A�nfvncc���!�)�]�����B����xf�Ũ)T#nGq��)�:zX�[Q��η��s���x^FFF� <�B�y�j�uc��^�����`�ߏ��u�W�X�S#E}��4G�>4feʧ]'=�����fv��q���2 �����r:�
�������@��2#�p9�W��C��@�wx�⏸ot�B9�ͣ��}�[�P����d�V?($1�Z��ʖR����p�ii��ܦ�2�g:��`�F,�ɪr�O�Rq��7�Z����9;(*� �5�-]ޑP��Pf��>"Pu�-4""BY [������8�TB���Y4��|h�֮���ܮ	��Šѭ�:z�ijiힽ���bfީ�mM���+�r��kK��T��A�y����J��zKo�R}�^^.��]�NS���O������F��*���f(�� ,��9f׿%<� �VXq��2.�M��^%F�-F�k��q� ܍K�t|���S���q=#ʉ5e����h�*����p�w�d[�-B�$	<���w�j��:�m_]cȟ�4uɱM1vhҘ:Ek������L5N��8�CqL뾄�ⓢ--�X%�`׻/ْ.���,�����S���`�ssj5���T3h����@_d��r1��'���/Z���Ũ�S��ܵ>��r������D3��]ŭd�����rp�n�S����"bg�h�U8ݮ�͒` �*/kl7 �_���7ٿ8N�����H|��:��Y��<p�E�h��Q�}���<�)O)����f���/��W�rpqz��芦|�f ��M�_�e#�s���0=p9�ec�4�<��H��}	C��nv�ck�@��;��8��- ����Ui: 3�|�hi5cLķuw�̓G�@xe��9 N3�H�.]���/���Y�?�H� ��p��Z�IEx�Z�0-?~��������a���i��1�?�D��WK�b�+7
[]{�f`N�����r2e��!�/��P�w�Ö'v8�5}[>tmt�V�i�ss(�x�N�|u���/�"5����#�u�N%��;���Ϝ����`iD;?�t�d������Rk{&U"����{���TP�k��[<����^������D����lJ����'Ų�Ϋ$�y
�U|�H�M���.V_�,B��.[H�s��X�l����g�6�����q�'��`aM���?U��ۊk߮<U7^ih�'�Ғ�0�p��_=R�kz���x�"��Qtn���ץ� r!̟M�[ګ�2�Cc����"z��������W�/ˌ"4o�ꗾ��]��&���k6겭�}�@��,�@��Sd�4��8�����m��zM�Ym2u����9����>��������Wer�Z�I�T��/�V�f��7i�C�-qdKf(m�j��0wf>���-�sಜQ)]w�.�Ħ����t{5�k_����Z��R��;�8�j{{Q�W}���a���ո����&{ٛ�`u>j��R��$����FX�����B�\9!O�?GW�V�g$�Ό%�oW�7�M����V&�_���P��A�窹�KWsf���K֤�p{�-�$
I��7����Pd��_�g^�J�\c���|ܒ��#�	'���+�B�0�}z\�*(D�m���nSg*�KǿMn�h��4t�����Z��yL>U����+�1�zx��uS�ZQ�!���Bq25�@!��v�>Fjj�� �5|L��mT���J�[O�' diҤxQN��\<�̙��E�G��q��������V�Ul���/y-�3���(Mk�Lq�M�G��yjx�s4�D�J���P^���@&�ңfF�މ~�s�����sJ�ǂ�mmtL��#�褠K�H���W�=����e�]�&$W_�����R&�ۑ���%�q�N(@z;&�`�3�[��n�3>��I���An�����VBԭ���S�#���j���}y�2���Ѭ}R�@;-_L��/���K�סg���{R&�?����DFW�p�����-r�E�5N7��'����\F�	���~cܒ妮�H:��k��s?�}�+1�<Y`��*�[��^�?0�X~i۲���)��>�]��������7�%h��r@��d����jbέΥ+G��[�o�_ q]���Cȁ�������!�QZ�pi�������Դe�Կ;u�+3�Wዑ}��ܥ�B�p����fmog��d��|���v���c!W�
��[��ǣ�"�Cy��ff�)������h����J�ϥ�#�[R)1)lpq8Gu)s-9v4 Y_��l�xj>p�Le�1���Ӽ(���EֆS�&��Xڵ�B(��kے<�e�cM�cw�X=<�5�S첤��Ի�bn�����O���l�)\���0ԨR�LگC���"�/) O�p_-���|�.aHnً]4�a�{�7x�D	�xb�܌���� �)��R��d�I궃R�B	��>PF��Z_^|3���������'*W�8e�h2�@����F�����te��/�{�}Ie�4eU�v��mll,3.��]fI֔�R�b\>ݭ��$x%ELJ��[-læ��+�HI�-���34�f����=S��Q5�QS��twN�sc���~tl�������7�N��4����N�u4���z������T�����^����;ȁM�`wc�k�m-�mx�&1�����Q����35����2���b���JA�� Cp[[*�T;|��4py;j_l�o}��b��B���e'�������)ug(y�l|o�[uOᩀ�[c,�rB�kn�/�O��i����%�G%j1�}������������L�%]�!9WB����5?_W͛���}ɺ���R2�;7����P�©�h��R��9�b����^ܤS��@�A��8�fi<,]����XNv�Y𝿐O)������P�	nA��LW��[�uF��ud��W����\p�"��� �G.'\�,&)3�ť�U��	O�隭�W3W|��!��q'�SiZj�0�d.��(Q@�J=X�+��lP���5�
\�u�#��ta�Tfwi(/��R����v�K8�b`�9�@�_��Y��z����E��������7�ٝ9Z=�m�bśT��#k�7��3V��XY}Y*�j,e�Rڏ�plC�����]����>���z���Pk�x��t::��b�ht�\_Q]	!���d��{Q^�����[O|^D��`����ތ��\<L�/��c�L�Zx���T5K��+#����Yg5�ð�F�&��=��.��%����וڛDb��]���9��6A!k[�KF�������aכc��[�q}��	=j��E"��aN˼+����y�D^��+J:��D"
��F6f�A�1�2��E�Ǻ%0`���FT�/��P&�]g�F-F
���fL+����}�����J���)��6B��ySݞ��,���*�0D�E�uԈ�r293���m)R���̠�3���>E}�H�N4ǘZY	w�����30C?����%�b��������i`���	;M~s�ŭ�g�Z�ϟ��4��Ͻ�_tp.ɿ���'���6vI�n��<�+��v�ߝ`��;�+�A�l�纇?�f�N	�K1+���;���q�^cZB�= ��k��Qʂ5*F�!km6>�t�\�Zy�6	���`��۾�����繐R��W&A��VT��2��w��c��b�2�m����ks#��wV��x�M��`�'Rja8e�@�W�����Ny�-xY����y8�,!�L��uj�8,'��uL��B>�^�Ⱥ�!�/�d��?����Ny�0,�5P���@��`P�������> }�=iǌ�uIS$RP�~Q�n�G��s$'�n<pxOE��R�$7�h�8��4Z5CV�Sjҍ����.���i��^�3�~�k�6k����Kͷ�y޸��@2WV�|��9�g���$
�s+��_%e��o͚�Te�
_����
�j_�Mzgm�>#"PwCn�=�|r���d���x�8�䳸K�A�=�oXVȊTn.R�(��~�lՙUd�/-��mYl:&Rlҙ�(=�*4H�#Q<�w��J�փVj�7�EQz��%$u=���]���Tn�U��Ў��������Z0���b��[[qLW��b���vB�<0�^��tUx��GX��������4T�@fm�%�)����ׯ7�z]����^}4Z`7�D�q"ı�;���@�q�E�2�p~\?cz3Y���w &��0vJ����EZ�Jy2?����6�}��K�F����Z]K����ʛ��638#�l��/ij7�c�כ�(��
'��V��q��G��t�m�̨���?����b��$Y��9>(�,k�����}>J�e01�/��w�V��3�֧Wߧ���-��;uɖd(�2�I!�N
{;Vq��%i::_#�⸲x�{���~�z]@
^�B��l���� VOB�nm�����l�ş�)�u�W>KG�
��)䭪����n-⤭>���
�B�~�
��#�B��E��A�������cXK����S��Myt�:I���*��|;�Ⱦ�~�P��5o�=3�_�<14���X�j�N�n�fӐ�8[ t�L���_r�3��b\
c�Vb-Z	�1'Q��J�x�d닕�־ZR)��C�u:H��/8 ��2x�Q�5w[�t3O;j���Lc۪�C�3�k��VW�+��C��X���ӂ�����G��F�͊n�O �[�q5��w㽉�%,D�س;�0�"D���S���ovt?�3��şj�e\��_�D�i�Z�#��e�����~��bR�k);�������{ G�!"ͥ��ovQ
h������Y6�	I�{�T��w"(�}ޑ�
I�b��a�[[`��@�����8�|�z�l���>A��XoԌd6'$��R��gx�bNp���[�q�Nh��<��A#��3�,��=��u�^t�yFY��40�S��Sq�렌��E&>�Ĥoԍjiűa"��'���Y�#�^^���uY����0������6�l�%or���y<�!�ln�n�,�gW+�m�n&Y~N�R�b*ێ��|�ہ+�<U��N;��)X!i!���_��Y� �$��&���.J~��n�+���]�ܿ1�cNx9+�D	܉�T���O�8������_��c��b�=����s�9��G1�����֣��JO�����3Z�P}'��Z�S}��cr��䁉�/l�o����t����Α+�mY�R����٧�����,��[�SG��+�R��[y�� l^��.uvypm]�x�A����{�?:���l"@~gI~ga����n�o�p=���*m˸��L*�������B�Y	\A<����8��"��^���\�0�_�8������I<�n��|'�I~k�L?�VQtron�1bK?GzX+��r��ÇP���^�!�ԝg��[��7���C��Ҷh%�ytE��te��qU��v]bRX�d��kv.���y�ܲ�s��cW�E?�</��!����ӊ�;�4G����u��nѼ��͆2��E�5y�N��ݪ��T��]���U5�����<9�CO��I�SYd8��^1��G;b<��zfk�fk��7���fY����F��g��r�zK��愓���+��'�.��,���,����Id����uu������D�(�B*���~FcF5[�h�-aΦHіԔx)���(NS��;�q�D �CS�aY�����;�esVO��L�`a��,�-ϝ;��2�a���a��i�ˆ�Mdӎ1���T��TL�O������9�9<��S�ɒ�降��q(��7������VZ�b��.�����y�= ��-�����bG��Q�6J��F�����L�=���R������X]���#1
5�z36܍���U�ny0�,��Ef� �����P8e6����,z���!A�+j�o>�e��C����B�̚�g��|�@m���^��������xL5ή��A2KN%�G�����d��EE����`�6�Ʈ��ў����z���E��%"�����:	̿�aeBE���E��X��S�b��:����EǱx?z9��P�O�E>�ϩBNƺy(mKN�l�#у����><�w
P�fU����,��[��77��ѯ�${u��)zM�F���Λ�e����U��G֞��=y��'qm�G��j�1|��ݠJ)ʃw��=�[AW���A��TU夂���[�.�eơ�}�zJ9�+mQN�Y�U�ם.e��O&G��ŭ�Q�4Yxܩ���L�V�K1)������I�����,��'8VF/2�!I�z�Y�����;L��`�L)b�D�w!�pH!'?u��'w�ɕ��-ɯ�yI���q�b����W�C�~��6�I���e5��z1��֕gq>���Ք�:�d$�7S��}s��2b��u�F�p=J���md{�LA �`7ZI�<(��� �H(z�E��j�����[dWQ�ѣ��$`�0NS)@��Z��`�ԕ�u{�6|.�ol�LI��JM"��-]�_�m�'����	���n[d `@8-�*����-���`ƶ6�pf��"`0�������?�7��є�sQ!y�+��KeOi�lr4��cX�3#���Kfs�j�tė��ڃ���z���&pO�r%�}�.���󐎽o"��<<P!qJx���[z�RS�^�U.f�'</f�oq�56Gu���\�R�nvN���_�7��a�q�������\��b�ݳ��L^9���ᩇ��~x���!�W�ttI\��?�z��6��/tO��TM�;���G�6�Y�ҳ�9
��D��O�����@��_	39�����%���%��7	V�?�_ �?��$����T�'�bމ@���%��7V��̂��(��������@��������+t}�IHHD��:�}�������:��0���:dc� ^����A[�g{C�+�n�T�����5�L8��r^m��*��.�DcV�OL/�K?'�z�l�?�3�yl�������5�����ݠ}����t����x��H�[+�*B�bT��ߑ�_t��N
	B\Sh��g)"�)����Z>Wd�4f���>�m�j����318zd'B�%��ܞ���W��-�vE�^�m����)���ĵ�L,�Z�30�W���U����[7����������P����е?E�Q�\q�_�ɑ#�j4�W 3��@����ϴ����9�Uֆc9e� ��;ۄO��c��v}�����Q���o���,kY�M>	?��`%;��y
P?��gg��x���(���7gnK7�t!�� l��J�=˔�VM׉�6�^�M�ߤcd�7���=�7����|GHdJf�p4)p���]�* �y'�V�'i������URQǎ+�U(�Wg���A[������9�}��y�v�c��g/��!����o>�m��㧍�$�k�kM�'n�m+l`&�E�=�e���o�1a�hi�
;��,��K�m�߷��+�ݤ-�P�_Q�\���W�AX�.������H46�x �{G�6�#����l��\��kS�~�[�� �m�q4�%��+��$����,ƙ�[�+�WW�=���g�-�r��A{�W�W��_ �24��ĹW:�����}�&赯�݊o�f��u�{����0��j�l���c�V�m�v�����ـ�7�e��B{{{�~����#(�l�o9x����ݰ����{FK����j_�҉�f�s���j�V!�J�wre��reӗt��f��3t���D|L���4����/�
��V���mJp GPh�� �y�����b���G�����cM�i�=� ,�`υ�F�hj"�B��?�V�ޮ�H��Č����Ə�)q�.��p�.�S?a~m_�S��\2���lZ".�/��=~�͗����9!�n��8œ��u��1ѯ��M,.�G���l�Udm�?��{�����oj���Ɔ�0aV��]aV�V��g�)�s#/1t��DG�yQ���`���F���Ƃ�y�� �֯�+�W�j��r>���@D�R�2���c�j�{�x��V��/�4T�bu��6l�JT�8��Bx�D<�F����1237?�^	���;�>��z`>�j�	�δY�4����5�m!Ci1��F�yЇ��V{�����6����p"�c/e}I����n�G��bݏ�V���z[ܯ�'�9l��7G��:r@�6�|���̇���\�&.�k�Q!_���rsm���؞VFdwyQ�lA'�qK��*�cam4�p2a����G��6���'M�ϙ���?:D�*n��g���ŗ��Ro��X_^
����xnO��Z�-"S��#��׬�r�zT���X�d�$�x�}�����KoS�,dm�����D�x��t�┬����D���1�7YK��GP�V ;�����vu�8v���$W�4b�� ���D�|�ul ��JN��4�͝�%��Vs��p�n���mZ��7I��ˀ��.�&̺��W���m��H�X���J\c9�0vH�MM���r����\���1ă��&�ܢ���ty,T}����ܥy�CWt�M�l{{�z0�zp¤!��u��CĤ�X>��b�`n<=�AB�ki�5}6�=u~�V�7�"�t�m�p����[���=e����&og�V��/�p�ז�3b��(��X�E�e�6�Jǔh��m|.hXr:U�HPml^�"n�B��I����X�`��N&6���,��_�޴�A����a�4r�.4�/���>��%�����L�|��5#ٺԶ��oG�d�EM��U{��������=&�?�y����/C1�ĿԶl�X��FY-�?��ŞjD���J.�=��g!��i4p�q�%堪�\�k�]b�#C�_��t鷓�>���*q'{����%#��^�j�p�ޞH	<z�/�8.����l9�'_�Q5��Q2l~ظ�ͰMS�Q����u�������F��C�6�������܇U� a=��O��͖Pf=fդY�>}?+C|�p��X��Y|�x����7bw�ׯw��K�.1���'�vUt�I��bTcUA���(�Bv�,��3Y]b���>Ԍ�x��Q���v]�a_}�q�p����U{��q|�ك��ǸMu.we�/�浜72̵��2k�'�&,y���v4��Z7De*�����b㔸�Ƹ%;lBq�P��ٵ�N#�O1K]/��vA<�)`<���G�L�8g
`oQ�:�?�p~�Qcx������Rx��M�cڪ��~��u2�y�O�|؝;� ���wF�u��<]�������s�7V2���a`e��U LL,6۸#��S�SSSV}��+�Y@���{p����ߛ
"u
��R����_��qȼ�^y3Qh��
�HNE'�w�þa��x7�R�B+%�bu1)��O8������b6��۞[�0��z)u�bOO����gb��HM�o�;����U4^%���8l0ף�g?��x�:��1K-�|{r�e)	�+op=n,	�yV�(�*�֍��Y�r���sz��7��Y��A�57����>�o�D�aм������֙Z^�%l�Ͻ!����t@J/�5s�R��݉]Qy�f!�j��)����G��楀�P�v��AT�c����]F�����*K�V[ .*�դ���'�k��b�~Rғ�Vpb�ˇ��kMV��4���ҿ`��WM��W���Ɵg�k*�]�=��43S�t��!�<f"�K�ؿB�V�7�X����o��6��Z������=D|�:d�%�_ߥ�Bm<c_p����ۚw܁@��3�@��~�ǟ�5��.I���$ޤ�D��R{����r	zx��J�z~���y�nLtKWjZ�Iu�2�G엣��,�E�1@:W�2�e�B�� �TZ���p}�t���I��;gk.��Z'�w��\tqG6�n>4������Y قș������#�1�~|:O�i: �U�c�A�!\���M���.sO��f�}q�&*v�� ���/�5Im��Ffl}�ٚ�_To��ӼR���'������\J�Y76��~�<��m}XʥC{5  ����mԤ�+����]�]�Ƶh�H2W���Pf&�I�g'a���"������-n���M�R��`� {����8�����Y@�Q�O�w.��x�$����7��ЉcK�S���	"�n�_g9C�F,���Aπ��G���0�'K�V���sA]���Pg!���4NG�>5q�L]��H��}�w+��>.Ԭ����xB���^�BW�U� J�U���h �ۆ~GI���8Z��P8�m�ץ�)E��G�ڞ5M�א���ęC�K/t_����Ԡ[��Nj�*�w[�aI^~�@��e�h�=�NMݲ�=�b�JϽ L�Q�3]�$d ����E�v���"��#���R׫�7�Dj� E"�������u)��Bw���Љ9ð1!�;�?��4to�a�����X��	H��]�փ>�µ�50�"�}��E.]9D�&��1Us��n�jІ�D�Xm��7��بǷ��[��7)M���D�Yl�.J?�a�q�ٯ�]H�����J�SV|������	sUe�(w�&N�^��j��1�g����ɪ|�wƛW�7g���i��1>�]��C���O:ޣ�R��*��P;�=&m�rn���0���w�p��#Zi`��.�ׂ�W��S�*�6���u��y2����ET����Ε�5DU�k�.�>��NdAI���wΉ���Q|�`�z������V>��1������M�Xlg�.��F���5#�X�N�H���ȓ��3�d�#�4�16�t�����n��U�����!��S˯Z��P���n
��(�+�߉��f�:�f5�\I���>d�*�Ib���Nׄ�����SY�TA~����0����̢f�l��NH�ӧ���v��H�q���TZ�w(�?�E�o�O,��tXo�ay"��aL"�?���9���!LO.Ht��Y&�|����M}W��p��T>�m{-e��ǥW�Dͯ����:镅C�����x0?���jML&J.7���cU����%���3�i���$_{�M3�M.���ۋ�|q��� MQS���M��x�k1������"ቡ�5~�G@���?8�JCB���6����%�.��A<��$Kh�^���y�ܼ�/��{���~���Cr6���v�w#�q����^瓜:K���]Ľ��	�����qM�sE<�u�?�j�Y�h��E�̷�n��%5�p�YnE^[n��3�����ƺC���O�!��-N������譡��a�f�"w��L�ݥ��,f���a�.����i"�-����l�������EK�ʃH��;u����N>}�F�B� ���jHX~���=y>�n>V���{ay���l,bMϢ�_���7dt��x��26ͧ^0pS 6��5�w:�g�c�(��kn��6)�x���3FFN�F濧����~�����"+�� ��]������e$�k���?��&�1����5Ɵ�:�7�*2����p_��QS���/h����Q��>U�b)�6ݶi�:�4��h��S�Rҕ`����бe���R�	�c6ӏ�z�o��gy���%��R^�+�А���♅�]��Į�.:3*l�H�ם���4��·�|>T���T�+QL]F���q<_}8EV;�]�b+0>ouqq/d+$6~�, �)�`I�@^��޳|�*l��v��d�`_��@\�sl�����WjeR�.���{I�(�%��V��N�BvB�̜c���C�v6���W�y8�C�?���#4����QO���2s)����k>c��Nԣ�%R��;���s���|o�֣��Ӆ�|5���gG!�������^%��*l�S^dɟIg�u���O�G՛#tN�.z��M��8���5��i����ό���y�ȥ�U��,>̀P�7�Ɵ$�[��n�
�0�*OM�5��r��ta���7�rZ��@W� ��Kw�z�DU�g�&�'���v5�Kd�E&= �! �dk��+]a��⏲�W�녇�t4�~���+�3��j�Vr��9�LC���Q�	)t��L����(K��T�w��/�Ԇl:͍sfҹe��E�WK{�BB7����*-���e&��'MԱO�ؚ��x�B��鉲��"�K�k������MK.=��p1���y�=����PH|hr�b,^��Ϲ�w��l�b�f6�<z�Oʽ��қB��$�Df�7�p/�|��s�;U�1���7h^��V4��?K㈿�������N�D�{��)�����_�5���o-_#O��SÕD�c�~hg�䢸�O���J��>��`���|z�� ,G6�iɵ����pa!,���P�LOJU6�������j��!�����&�,Dw�`�N�YE��W���w	�d���'j7oa���0A.�coKl�����b��[^qtc�k�@��LM��'�o���P��	�;���Gl:`����(I�e@)(O�]iB �q�W�>���K%�*�6t�~]��k�ub� ��;�����N|:�침��{�oU����'<q�$�T>�����ys��N�R
!}4��-t���Ѵ�
h�?�e6g��Z���ӫ�g1[���.B�B1��3|UFf#Dڋ�by<�K��B�?�W���3����d�M�����3a�	~�o�!w xh;�na��Ĵ��A�Q���)%�#W�`&Uǿn&�D��������MvN�R�U���G���Ն{��9!!K3�Wϟ��8�~̲{B^`}���j�k�d��>��R��?���y��Y%>Xq���pGy�j��I'S��Cg�*��D�k��=ZP7���L��\�^m��p��UH�%>D����$�������<~���#t,��U������M�	�$�B%�7L�p�5�����J_=pz�� 0����/��iĊ�W�v^R���,�nt+�A�Y����-�%��g���-�x��vt4z����[�~�����Z٘���2 E�*ݴ���o����L3�M�*J�և�ɠ��R�8�9Z���� ����Ak�����P_{Io�^	>�v�p'X�����������]n���m�L]�̤Ȭ�!�(SfJ����1��2���)���2Oq8���1��]�v?���=���Z��z=_�����k�j:\Tأ^/v����uE����R� }G^+il��>ɀ-,��su�nl���R�ŏO;+�[��[ ��D4�������s�8z{-8賡a�/�>���~
x��$?�7
NF�rg�m�B6�=�iz���Ʃ�����眵�KtZ
���:E����O5=�dm'(p]*�H���B����ss�V��E�9��>H�A�H_x���I�s�}�m�Sfqc6��/o����C�p���J�u�����=���/8[�_��-���P`>�iKp���ε"�y���`6!���e|J{z�ʂ��p�ιy~a /!]���7�[�c"e�/6���(���?����Ǩļ$��-��+2DL�u3P�
ޡ�/Q���z@Cu�V�iH��8�P�{X$Tۮ��?uj��^ps��[WDO^*��nN����%��C�gdt�g"��/��xC��E��%��B��S����ŵ�z$C�b����0eu�9��\t<����5�=g2���+�5�/��3��e�9['a5�G9���7�뀩��.ǧ �O��]2�هac���8h<��8��腂-{���.�=6%r�oo*��"�2;�C���E�J���Yl��6
K&�;`�=���f�4�9kE�=��}��>�rO���}�<���	�R�{AD��e%�H\fy"��ۄw�f�i
�E�梔�tv=���~����}�zd�^�i��}<d�5��kg��Q��j�=�{�P���0�6�1��lW� ����BH�3�����f�Z�>���s�%��\	�Ǖ�LOd��ٞ���p�{J|ieI���5p��Ԋג�UU"�:F#�n��쑛��[?��'� X�**�p�O잷m�z�lA�k5�D/
T�/J$�+(�P�J��Zy��'_v�fХg
�cQp�^챙"�^{]��4Z{IDi�t�{�^����uD�v;����K he��B��k�(3��O���}�Xk�[�wZ0�(���[N���t��9����4?WT�x�7��E3��)�tW�_^�$-~/�����U@;B8�����ʵيhx܊����,�kU�������mω��, g~��lf��"Ҹw ���,l�QT
�$z�~��r�.$P^ ����߼��U�C��\��ֿe�0ف��?��d:���&�m�`2hǯ`*�⬿oL�!ꣲ�u����R�ZC�ݲU�v��Ր���@�\b8c�
��F�}�� �2�q"� `gO���$�y�#��y�=����q����:�8g�`�t�.t��B
Ȋ��S��4}�F1���6����HK�ٽ(W��W��c�)����n\�iȗq۬��ת���.�x��g(7���?./=o���b��)�y���R�bL�	�ѡn�۟���kfC�~�'��S#��p+Ng��Õ}���z�I9��?��^��U�2�m���1P���=Z�a�l�	�:��>�Qt_�G����P_��[�Z:��ON���qe��G�p�^ n���\�9R�]Gmi�V�ȯ.+�ߡ�������V��
@ș�w~񫋂�5�����{�G3���c���{���V��/WdB���wVQ����"�h ǭ[Ğ�zY���(�u8S">E(n[fɷ���Gr���B���aZ)H�N+6r�R:"�e�F� �W	u�Q����S�6�V_H�?j�|��{V-(N����(��:�|�\w0��Z}]ۺ�{����#�a��ur���z�	��W��4�7�)�4��B� \j�Wj��7^������J�θ�<�7���x���p���V�>���.?��u�
G�2놧��!��;��C���+�ƕt�3ٝ]���
ؒMk�3�_�M����)pq���Z��E�U�{	ɑ����Ķ)����dm5��h�-Lz_L��b�(���/N+��+f؂V<J����t��u��@/9j�DWg�����%&��D4�w���V����t�1�l����A�ج]���S� C��)���(�bUT0:�?�
@[��+�8���e��3uG��u�6t=�_���N@��^?V2�PI/!�v��0hX���솘��<��>gJ$��h�����eFھ�%!�G�&��R��/嬝�C��O��4/|G#m����i�&�f�D��^o�=�A��ske�c9�Iolǣx���{jq�=���9o��\�����'�,l|%��� �[�@��$y�������L��E[c�L	�;W{Z1䱃H���3DM��i4��1(�G�bhf��
��x��x�� \'s� ���G��Y�D�H5����G���Wq��#���"�#їP_�d����7� �d��X��:�~t���p���E\�ФsxFF}th�$8���7��7�e��:�Yw�� ������f`�&	�˷;`o2OF��X��� -��8�}�$)���O*�H@��HM�Ϙ�J��Ģ�w ��:[f��E�����^�HU�z��0����9B1�S�T�#LLv�{�U�lRT�#$�(7}�u+���C��N�Խ��B�b0]��JC~�M�C޺��t���Ǫ�[�#㵊��ď�3�(����S�ſ��eS`F�hҹ"����e�Ѽp������(
���	W�*1��v�`�gR�X�������?��� z���gT���L?֘��T��m��B۞��v���9G��]읠�5dzFd���`�������͚@[QB�g������A���M�a�#��"!�P@���ܜI��dQ\x�F��.�f�dC�J��P����]��
�m�����������;�.���iq�yQf���15@5[c�rqT�hх˙��J��c���t]����M��w��>���\�-� ����~��n���`���E\�*S *^�6��-���:u�L'X$)�ג����}�K�q�;/���/�
��"<�yzgBbz{�=S�E��itz�[���V1�r�U�2�7�1��:�΋`�P��b9;��[��Q�<�Z^��9M�vu\]�:���W2�]5U�i����t�������	�؃P���)<��`ke�m yF�K�s �_�멿�\�c�t�n����)��vE��??��`�ǵ���ygi<^M����;�~7��)�%���9&��MpI��,ՃH0���gw�:����'��ǟ��S5,���sTM'�61�-D���q��Rcop��kQ�
FwzT0=!�v:'y{$����Դ��w�=��V��ơE�����^����_��U�c�*e�m	-ά��D����m�TI�cO�����n�	ܿ|�ǂ�b��q��s���l�ڴ�Z��q_��EH�.O&����v���w�4��7Z
f��D�l�#/���}N�ٮ�U�:����=9���-H� ��V&��_L�l74�����d;� ן�+\�5�9�]�¢��\�b��F�\�-U�1w�	��aDlʚ[��Ƿ|d*��i�����V�8��\'���y39~�@#�'fz�a��@� �aH��J��M���7��M2{���-\��70�����=������,�3I��nR7�I,�,zn|
�Pe�����/��:��ͧ{�VzI[Qwn�jG�Ʌ ����J]�"]��T���I��7�+<��(1D��\�D+�NG4�L�%^�o0U:�����P�������E���3�otB���@�9� �B(��жD?U��õ��`�gD��o#�d����0v\21����s�d3�����X+�QI;k8Bޜ&����ǳ����e��y�����Ƙ���vXl����E9���6�����va��7�=��2�Bv��Tߺ���/k��\(�����%�6)�u&���{{cv޿�P��x�o�_�(I��r��??Pz�[Nse��a���^��7��3|N�<� �g���!Iey�j��w�B�'Bb����ph��+�Nx@2�����,T����f`�����â�\��|8��JKi��n5qä���i���UT�CEa��4�]"lP��K��V��&S���r�����AY���7��I���	�1��)�|
K�����3�an�>��2��h�3���#�'!^��U���ij(��E��;�Laz�"ӳ��BQ�]���A�)5�L�s��T�Ls1	����m�%˘�N#����g����4~���(+8_t�V�\:uL�|2>�=�3��	ix��K���qm̔آK��;8)r��3�ͽ�M�~�\�'xF�̤E��A�+7�L��kU��sʠ�V�ߎ���{ul_,�]q 7�\�E�hZ�T^f߮���ʩ&��E�^�,�ߴ���S�f�ה�������>$�n���qgS�l�-��g����N|�}Șk߶�V�DsE�����*Ԫ���?2/�;��K��U��\jy��'U3��/o�o������:�&��R�\�RK���Mö�k�8�v����H�� ?T(rf����wiwU���[�TF�И&�9U����	*�����d�Qg�DXP���h�����DC͚���:te����3�ߓ���:v���󫮮�l�ט���:ԕ��u���8-�qӦ��@�4].��f|NĦ�*s8��Iz����:F��xDԔ�6���hb�$��5�9�P��b<e.�@��E�[uf4�*0
���s���i�(d|�w)�M�dwM2���W@)���?�#�e�ܭ��[�)6j���ޑ��a�rc��O�[uf������K�D޲ �e�}�ũwʫY�����!w.��teb�_mX�� Mb���W4�5�9"��֝gl]iۑ� ���A�)�^>G��Z��T6`� �zz���k��xv���Y�(�I<��d�fd�P6P�Qk�2/�y7%����:�:]��Q���ȹ��R_Q>�z�Ӱ�N�~�wJ��s�ߍwDT�6h[\���I��ҹɎ�r���m�ŖE���v���;�T)�X]S�]���vc����#6Jr��dȼ`u���G�j�gq�	�s�|�C���.ՓB��NS�EYt�IQ��!���K����q�(��W�s���I����7�j�7����������t���	�^���7��Ê��}�pG���)�X,w�$�����r�^Lt�pd��\�����ƙ��9$����̩�+�U����j�UD�x�0d��XU��g8Ը�0�����[ID�PL;�_G�#E��sS�bь�A����X����Sv� ]�����v~����wV1ErHk^���n����đyCMowJ7ݠdr�I���Y��§��Fwg�W$�jU�=��dJ��{C�4���}NQ�'�����i��ɚ�}�7����A�3K3p���e�L��c�_��z�0��UDG�ot�R�+q�f��$�~�T�����^0֒��g�A����rs�m��߱��w�����3{�
,n����P�"��L�l����>��t
qW���w�,Q��K"���Esi�h0�	EKE��p���韓��z
T��7��g�ly&Ip0v�_��Z�Q�jqn�7/± �9;����܆�O�[��K��&RHA%�wy�1���l�}�O0k_��'΋-���uE(��T����H3h�|�1#���ct�|˹N=&xփ\R4(�=��1�1@�())�P�gn���մY��0²��cPl�Fz�Q�v��}�fp���3�jȷ�+���7��l��f:N>ʭ�-#�HK٨[����?��a �WO�U�^���-~��w4	,[��&�>� .�P
㩅���L�����嶫T�T0��*K e}V[���"a�5;KjP��d FW���㒊����ʊ�Y�}� {�㻼$��(n�lw���%��C��c�ؠ\��p�h[^I욹HA�����R@�G���3��Ӏ�$�����okdP_x������ۊ�	�uF����ϩH��X�(���3.��sUvQvxq5K ?1Q�+�{I*����Gs���ec1��74���.�������^�MB��A��1�G���RI���ސ�َ݂�J$a�ݸ}C��~iT�͙��u_�Aش�hʆ��>XpndxRu2}��0�Z:��y�����L���Bx����z��*������#Ώ�F� fB��N����_����R�S[��J�DP�+�C�|c�!}wBz�']�zPV~_���K�:�AeX����*��}���?�+OIQ��=p*��
���Ƃ�f�B;P�k�����ϝ�����Ef�~e!��e���7
�������:���I���=*?5��ͻ��t'�#4���B
�go�l�>/*	G;���,y*�����ցf�7�[�� ��j=J�%V�b�=��ѧ�J�v3��1�7܀37H�Y���ɱ|���**8%%e���|9�[3PBd�spi�N������p�|@^cb���4&�36����Ow��磑V�&��4_T�L-���w��|u��&��~�h��^���UZz@�~'\,Ze�7/�^: �"!w���ja��ĲE��'^�����Ra�h��d�qʫ�1=�S��B*;9w&>����-�7�x������=xAv�l�3�_�א��:ǻ��X[��P�%LYǃ������r��Ie�������=��VlA��2���K����Q�M7����0�DWg��<��Qc��S�!�Y�߲��I�Y2���h+g�6�����E"���}�|Co]���"\l���l�5�����*�8A��gM�1����2G���_M�lp/�_�F��`�;�uU���~3�V%?��� ��dJ��6���c�N��n�ڜǣP�>��_��CD�n��-e^�tʹɠ�h���dĝ��גܖ>�#W��6����M�����FQ���_�ꮕ�M
�?|���� ����T�u��=s���|`�چ��V��v�������3�p2��W���V�$�Uy�E{�����l:�<��*Ɛ���(�A.~��WB��A�5j}ghY�~�1.���+�T_L��Z�l�O��خ�<��|�*BW݉�ο6e�8+-	R9pXy=�0��:������b�.[�OJ�脤zc��6����G���qB]�UNf�o��M���Ԑ�;6M������y!����$Ѝ�`�)%��5�a�?�:t���1�ѣ�I�q�#3�?�H�j�Ϫ����j�9���������ysq�5����aD\$��#��ɕh�V�.t�'�Y~�;R���S����c��T�r�P��{]s��������٧>"�?��|��v�ˡU+���n�Cԕ''���8ɁS�3A '�����d�c�P�A�s*���sm4U�V��K#��N������%w��:)L0F�oа4���F�Z��
P���L�U�M��s��ѓ#�O(�g26�6]&N0��I��5���?�!��6'?�nQ-�:,D���+��L_�X��VS��_���C�5E �؅B
��6�a�	�M7�McY7ak�Y�P���X�mˉ��K���%2vë��Нxi�0ߠ�|*_��(W�b�nm֦T�)�7�_Z��W"���x�D߁�,{=�H��?W|V�e��.'�=��y������YtuM\���/��r��Z�E�!�у��>�h�[�5��j3o�:ڋR�O"�l�uoZ���7��g&�rq¸!��|������Y�m����z��������omN7{Sk�r/�*T�r~�*+�J��?�~CW��������P�ʲo�Jw6�ɡԭGrzU�OH���/�M�h8����wL^�������V�^W��=�i�Q�g�q�7����h�՘EI���_��FN�L�^v}�J� ��%t ��a�aY�%-򦶬~��d4C�����x��5o��2Mϛ��Gf|V�M��������+�Z}|�}�����h���>��@��^�C���j���H/a�����<�#��S����m"S�)L�T��3�2O���A��;����rUUmЇ�*�F�/&�P��)TU��<n+:,���>�����Hj�1l��*>p�ĄD��ۚl=�q��2��K�-�y�E0���R�i�Hg ��>՞b�Y�ﶫ���iv��՝��\ѿ΄�Za��,#l >tt�g�̓�zXm�^����f�O����`O��z��A�R_o*�")Q��K��_VD`7�wO�����⎴��j����r�7|�Te��Ff�$�{�7E�X��s��I��ZuKҿ���Ę�.vb��T����:s���#W5[��ݔe�g�81�s������K�K�_�\�%$/jH�O��nΙf.��v�U+�N�����k_�,�]������U�k��/�c|VS|V}}��.�{v�rn�蚬zJ�f��5��԰��";�_	Z�>�H���n�b�<�;|*NӲ��1���@��L�RA�e�a���EjY6V	V�/:�G��*�"g�N���[�W����od��7�:���MI^`q��ԗo@��։M�5
km����2��0P̺
@�IZ0̶���>��l5A�U6����f�<g�8��t����M3s��ZԢ��6%ډ���ʜ���ֶf�����h-ee��/1���_K�vF�8�g����qڝY�p'�zWI5@� zR��eM�K>�T��P��t\��n�sz����%ܿ6����c���i���fO��q�������Ykn<I��@]��m���O�5u��A��Nrb�9��o�e�\t�Zm�x��u��Q!P��][bӃ��ٽ�\��2C��K��J�2;�./�	�f��+�,/[e�,[u���5k?�
��s�}6v$�|*�q��8��^jz�:��=��2���s���k���~�e_���yp�ҷ:��|�tb>�q'@?�NPp��-������T��h�	�g��K���y^P�D2F�}@p-�jOK��Fv������e��g�-]\U`��F��D8�<�1���z��v���u�̢hw^��M�B���:�i��y�-~/,B� ����L��Xޣ�~oc&:����q�s?ێ�q�h�8[ad�"�Cp
D#��x���d�H9�ʮ{�>W2�5���i���^��|
�/�
ְ8=��Kt�v�:rd߆O0|������W�:��#�AC� �tqG׿Q��g-"'[�����긵o�)����:y��S������ ��ܯ��������兼2��m�u�&B��D�$փ2F����!N&�qA����#�K�G����?V�j:���
�:��I�w�����Ȭ�b]0��>��M��??�̥����1��������R���c0ు���m�?����M8�8�ghlE�_�Ə�� AO��z��h�A���O���S�l�H�\��r���4�Cj�B�8�N�с�d\i��4��駔��&�RPo/e��t�XJH��Z,.��8�ԸË���SD7$v�L���X~&�8[N���s̛�#��s��p"�����8���<�FDD��Aj����g˼�saJ[_>�\8�Dj�Ճ�?~������������J$
���NV��w�?���*�(�äƛ7��;(p�?�'����]��W��]�4����U�p�Pp���^�^����ܿt����m]].�C��H�Qؚ��S�;���FH��.!�cpP�Р|)���t�
�gg�$]��K�Ŏ@�H�s@qʡ8�`	YW����5D���۝��ѕ��Α����B��N��O%��N.�445Uon�Ʋ�Щ�$4�������ǅv_��+.C�T�zA)6<��uu�5�ޢ��fU�]$��􋋋ٰ?SCH�� �+��P�/��W�9`��LS~!]���	P"p����k��-#=D�nz��ťW��5��� \܄�.�@6I�1��Z}�����Hc�2{2�WZW3��& � 1P	1J|�j�C�u[�;��@����]3�}��@��M`��o��ӝ�3M�D�C0�Ll��B�|����a��e3`��P�+�d�I��F�9����Sky�h�_�VG�J�b@�6���P|�0�Q9|�:a��]xZ�@H���}�7H���cmm�,BY=1�}o�9��ty�H$�;w���{+dI�Gi��m]������5��+���p^H��e��2b��쬬?DIm��-�t�=,j�f�J`6Ε�iݓ��b���\m����)+�����G�¿a�x��/��vBӄ�B��TPXHOj�V��=��ÇH)6���M����+ߺ�{��Sg�X*2��c:���jj��K�yS��Ǐ��_�jY���j1l�B4��n��ul�^�����4:������G
����}а��|�m�+?�]�?0���XtJ���3R���+��Gܿ)�hhj�K��(��3�3m�=@0i�jbb�+�A�O=Gy`�
�!��Qb\|�bG������O�<����
I�3}��
�"w�<�G�m�:l��>^��T��펙�|���&W��ɾXۏA[2��h4��RM�3^��\b�M�W��8�}����	��[�����<�Y/)$o0	��p�S�2�pLj(@F��$�l��Ҧ:v,���6��klj
��ӛoc����q�%C����BA�*���~On]x��YZ�~�f��i{���^�vs� ���h�&T�0�����w�=|��C�Q�iM�W��?2}�O2W�X^�G���������R?@�W�Y~5���Zd�PAMԑ���9�}?�h-�}cEk`������BC\{�Y���֩n]�A� ujr��Y�,oƴy�aIMZ�k
�Tq,{�P�	�+~+нl���l�(�����l�9��I��|$�w�@r9��m�_'�ꨧ3YW��<J���+����=]�}}��F���~�����a��	�\8z&&�ngN�N�)P3힚-���*�����ع����8�-�F-�빜Ej��6w�nі%�.
q^ӽ��������:����T �8f	�
[n�+���(���d<��m���K�����-�{X3f�82����T�[W��\�|��5�t��3�6���D5�_Yzz�������h�*�-5�8Ja��t%))I��Iz�W��o�ځ��{����S`d�>N�(U+M.��~|��U��Dr75y�P��!w�=G3�>6��Dl����}�cg$ �o;Ȭ�o}9[U�ƍ�-�#-��$�Mhp��:4�e{�	:7��'�(?��܄��%�E͊ڏ?��2�p�բ�<�9ML����F��^6��c"}|���RS^ZX�j��~A�b���J#F���l�qUS�O�mll4p~����� ua͕��s7��m���%����q�HY���3�ֿt瘛8����+X�>U��E״����g�j�A[��]䞣�[����y��`��V��H�C�i��A��#,F���z��W�,J�F�����Ề��:k��7n�8WfY�]�6}e{444t�������ޮ�q�aS�� �N/��.����ȷ�n��6��{l���3R�x�,h��u�P�Y����4��M�g��w���˿+��q��G"�^I����٘��c�^�)��f���A���P�R�hS�8��Ӈ�
�|1�ف�����1i�ò	6���=�Q��{�p�&���T���� +���F���l�L[��q��=w�v����ʰ֘�^^>�j8�=sʚ楯�oW�����~��`7���P���p.j�IF�(�<�z:�f��?TU�2^��K'+��<���e��Aq�����ZXI����{�(�~��_M���o��q�t�W"R�д�G��r���P�.)}� O���j	8��gce�WP0�X]Sc��\D�uez�&DI���fH�F��ٗQQ�e��|׆�Qt��?�c��8P���C�jum�H_6;7׾�H�ҥ���rM��R��!8���W��H��(�����ӞNߎU��)��*����O�	dڨϧ98n�G�Ke�`��1����� |X�F�yHH@�Vm$y����9pBd�o�)(!���s�y�x4��zxH�ٞ�C�)����"�	l헮W�����8͕X�i��c�U�%���(��h�9=��]������	�y*�6S�|d&�����A��A.���WD���?)�}�?��\'*����=�:�-wnR��ǟ�J����$>�= �v`���A@�+�)b��X䈷�wɫ��
7//�G�<||��zy����if���x��M�%,I3�b%����ͬE>Y%���Z��/(C��pۚ2
J�q�BWl�n��&�:�>a�Ɍe�i��9�}���� �r@���
����gzŁ��LR�VV�|��:LWA�*�v/�j0�+���Nc����8�o���r�S����qP�ִ��e�"��և~}�p�ɩ0�$�)�� V%�*)�
�+b�DV�HRt��	�g
��&�؁|$� .�E<��
pi�(�D3O7���..&�N6�X��<m�z^��׍vUi&�U��Sˬ���AQ���r���l�`��Fڗ@�O�
��,g���l2����
��9�*�j�IM`W�+�w#+���{��L43U��w7*�%��V�dYq���� 0���Y���p�豞�)�i11q#H��3���[W�2ɓxPR��s����S�{j�n��j�Ν����1W���	�q�	b�п{E��{�;�i�$���t3��[��Fku�Ť
N��H���٨`�uܸko���>�9E�)���A&�I,-�`
�z���r�>(��2�Eث
����rF�XܗZcx2E�cʛ_Y�� �6��5U�QZ΢�
����Z�,�:��p���i�p�:��$�W�����H�u�LYm/��1�4��+fH��6QP ���2�\[��hXP:ʛr��[f�&i�-�����*��Gq��.i�B���(Y��O-6K�x��{v�F���j
��]��g�Μy����4�7xFd���?((<о��z�ʝ�Ov�8=2����Y<�s��q��@�4s2��6~�+0;�Ñ��}JO�"��:��@a϶�5���er�.+�qG����\����é
\�������"��G4R�t��ߺJU\��Q����";'�7��]!		Ɛ��#"�7D�O �O�c6n3T��b�kmW�þ����ʩ�X��n��nsq��A����{Dr�YUa, (H!Ow�>`u�^����w�d(wA� G�{��;�Z[[i�͒ѮI4�^=+��Z+-�{`�.�;o�B��+�azh_�h6��jO�CQ77�z���_(4�ū��;7g����� �T�t8e�<H�]@��q�Cũ�����fgg6�/J�,jkk�w��1��ǯQJӃ�4�D>�7��eh���%b��o�h�RK���t����"[��E�VZf�R��CUu��c:S���ty�]�e6L�U��R�jM��`ߊ��ȈM��/4�Ȗy��V�W���%|	�e�)+�	F�L���E��E1M����Sy��l9ŵ�+ֿ8��8�b�%`���O��4E����^��������0���� ��:���͕(�U�^�ZO�.eRv���p���T8��#eU�r�aאpK�\a�3x�S���,�)�;4���$�:�ye�����i�#���߹����HQv�u[���~�����=�<|\��g�c�E�P��,���R$�4g��V.l���1����G��F��{�O� >J'}��W A8<�L�z6�Zr#�Y]�_��s-�4׿���������֜�?��J%G���{P��E[ME (�Z�G�Ib��c�^ށ}�,
К���ͷ�B��\�Ə�r� �fcc���oS���ވB����eC��� ���*��4Ѫ��+ߵ�Le#;lq�6P��48�HhӁ��i� �cy������Cp���h:���7�(W��?J �1�;V��Yafd��(jQ:�e��x[N@�,�k?����s5ˍ�pC��i!�w  �Y��tog�(�I���>lS���&����l��
����V����2K{����C
�_�x�m�4777����<q��ի�S}���Ĩ=�O��:�)Ж^�>�_&��)6�RSTV��-9O��y�}���|)��h'��4;�w�@�v�[3&�&&q��8��Lh�u1��-��-����n5)4��𭷀+=�/�*
N�j���:�Jԕ�L�#����5�B�_���n���N%����Eח��th�o���YҦ5AmM5�d�\�{B�E�kK��90�9��B'�&���#u���ᗫ��Wb�j���B�Cň��R�C��SU�w�.�'�d��M��TWWGv&3���f1M��$%�,.�QPQ���#3��^�Z�����R2^W$���o�|AEIa¬�v>VEC�b1��q^]�Y$\;p����Oh]9]��m����6��f׸����e��8&u|��H�9ݛ���y'7�#UF1��Zb�P?���a�����=w�Azjs]�J�ͪ}�n��e�%:ZQV-����:ʜ�cQ$�a�]7٨f�X����!�ta�Gh��lfJ���;�cVf�{�.��
򱕯:N;�ִ��ǉ�`���Դ�J�AL�u�̄nkC2i��Hh�[w{��H� ��D<s���n�s���չ���w�ٿ�s�\F�ž|�`�@�q}4*6��k/̀ei#����!�K�0��`�h�v$%$6�>x���0�e�#˽nRB��^Ʒ��ȐI�"�i�8��@:w�e����\z�<ϻM�#�v�`��+�����ߡ\�s%�J�VT|^��Y���\YZZ�V����XU�\�qD��ɌW(5�Su�y��	��BC��|p��[>VC�x����N��:���:1QzH����Cޑ�bA)���ߗ�m���d�qN��#�:h�����=yi�#� *,b�qo�]�B���n�S���'�Ѕ������|J؆)C{�_Ft��� �8��ɺٹ��?w�9腾�a��`�%�Ӗ��o�Ҥ_�QW�ENW^��b�gPC�)t �i�~�H����x�X0rmm�#S��W�,�VP���@���S�"�,i�� �X��K�Q��8�n܈<�_G�.��l{��V��J�I���Ev����
��;m�o�x_)�\��B�e��_���3b���נ�Os4��?;{J_�r�!��N�7�_�X����j�D��;�T�rF3+#��*u�CHfj����eي0���y'�>j(��3���g(ՔG�x.����*QRTʑ�s����"�a��H���Z�(�-�G���lT��Z�wq-�U<�%���b�����/i�\ G��`�����>z7D�t�`%�E����w��O�}}�c@�j�?�ܗ��{�i�|g�'�UG�dRKT�{�+B̏�өl�B<��6����9��y������sǊ �k=�@�5�2C���b�d�����rٗ��)����S�퀌=�>NN���7�d0����/aAĝꩩ�rgL��(pg�;��%ќz}J7A����o��V�y+s�`��[��B���������Z��Q�J3�Y� KY���3_f�E~_k�N�uԄ��^�$�n�(��V1��8�� ,�2��bp�������w�y@��+J(�9�T2�gjb��ȩ�嚯���@�%z*V�}�H�q��C�HSP())�7�N�d8�
��}�@�b�T���P\(wgY'����Z}Lg����;���w|_�+������C�6;?�q�?j���P�q��[T�	���&Ȃ�Z][�<�U�C���;&��^a<uVP A�q� �u�;&��B���m�X!5ԹW���E�1��~�HGg��Gw	VL��~��Z���|^^�$�s�Wy�����`�)��e�^k�C��H�B@:�|G B�\���l��q:@�uj%�w�w�--e�3�:�\�1%�w�w��tO�2V�b�Nþ�'�b� -�g��x5�"�9`����*�z���tck��a��۲EZ����H�\~A�	�ls������L�� ��GHx���]RXDď4ekck[Q�x�laZ8::�h~)q��b�@��H=��� x&�,8�����1���$E<I;��S3MK����:5݌9��Z<���鮾����,.˓�<,�W>T�ih��7
	��V�s�_V6f�j�BxhCz�n�bj���h]���KNƒ���Fl���i[pmJ��p~M͜�EU==�
�)(�a��g 8�Z����"��EG-
���d�֘��N�
p�윜��ME�C�/F���2S����+���)��yצū�7�|����uH5�-��KIm�-��!�]����za}k��<��V1�S;��6��r��Ba|�.e���o߶U-fv8l�4K��</�_�P�) ����]���#d��hJJJ�H.hN+��ut|�uu-�V�E-��82u#l���jzzt�5<���M�Q��Y,��7l�or��XR����cu��ϊ��P�{�
 'LĿ�8A���VZ0By�t�j1����y��������ԗ؞h�'��{Z�B�O�W����"�ʥ��8:9��&�A�t'ڦ�_�VZT@;�&�O�S����q+q��3��Y&h�Bu�u��08`s�k=��e�^�ٿf$�r�!hU�7o����TVAlZ��⌄�	ق� ���jRqFd��)Q֘���������׬�uR��dJ�/X�"3�QI�Cn�6t"m
�H���� $��q�S�אs�R:�_hNPT�a��Q/9GV�)P��J����/����8�ֈ}�:iNCM�6�r�JM�{sT��m�v~~���	�):�}'�}VRS=F���F��A�$�Du)��HSs�8��� ���[�z������&�/��10gN. c�]�����1?"�)3K�(U^�Q@x$^K]%	K�KjF���H�8y��@���ylՙя�pE�CȎ�O�l��T#Yt!d�d�~|�7��4�R?:#�y��ǐ�,v���X�aY�Yǒخ�ޒ^{N(�1L�w/'�"�g�������"���o����I����ooo#����B'F� ~�UgQ���	{�"���,���vG�]���%�&f����RX�d7e�%/���i�Gδ
�O,���Ǩ�H�����>��6�V�a0�)P��L�˿X� .vgx�u�6ۜܟ���l�����?PK   JrX�Rr5�  5 /   images/1c16f167-bc9c-409e-bb79-de4c62b914f3.png�gXSY�6@���c!��cE&�;l���ҕ�*EzO�(�t,�����
J�*5Ajh	5��Cq�yH��~|��o�./=g��ֺ�{����g�_����)�	����9}Bc��`�>q������ ��f��W]`0�S�o���a�=�3'�/yƎ�pe�00ٿ�ڴ��E�=��͏;����1SV6�[��`���9��w~�K�*�%�6׈�Ǚ#Q#�˿�Mi~?���u�Y}��!�+�~"|P���%�1[�ߊ{��}�z�|�/�?�X�~W�@z�3f����jC�?m����q�9���?h�lĻ�;x{/��YBS�"f�uF����C�<���p_�y'7|ÝWj��x���3M��#t�R��s����W&�j�0�pKb`��/{\y�T������;�g^u/��*Z�~��n��M��JH �h{�;*"�t9d
9\�fMϚ�ċ��#��.�]'o�&&E�F���MܓꝨ������8�➣�ϟ��X�g>�1��W"b�������9��p��ut"���xx�+w���ȳ��!S�|��r,�����ʫ��Fp&���B���R���!F�$�}��K���!��N�����ӷ�U�$^f*�=;�	��n�X�w��r�ܟ�@ԅ�kW��O�ީA9���D'ԋ/����W�}�H]���ǉ�3�P"n���t��j8��ܕ�l���eȔ�ћ����=��L�6b�E�h%9���Þ��3w{������1�I-�v��,?�+&Fp�g��؊z
?|��AT���{v���!�*%����زkAf��ΛsK�f��*���-��O=�BRO���'�^�Iy�y��_�1K�/�6����`nkk��1�	���Έ�8��8		��U$�1�hk��v6�M���9׆�<TI�歈4���ѹnNZRQQ�v��V�k}�T�ӥ����،����y��+��:B�JO4�4d
]\PX~m��v���ޗ�W<2w��@ʯ��E�3tJ]b��3 <BnDv�L���QVA�*?��mV��oߜ�ܤ��7iL֗��bV�������O>�A� ����ۋg�����C(�����[�I-���
�a��=[��������=FVfO������l�R�e�F����2�^l|��W��\ �N��KOx+��M|�������C�Z��n�G�������-9�C`>�:ឰ[��q�a #;�233���C�s+��0���?��M�^�VV�ec�>��
)��sޥBR��.���8�Ԥ;�����魶y�9hu����<���=)�r}�ֆL��J���M�ܹ���3�����|)����3!�1�Qi&3#cpk���C�,B��`��!Khǫ�W��\�|�}=D'D���~�i���R2�H�r��"�Qc��D ��W)Y��O	�8O��$�8Drqq:C`P>싄T��c� �H���C���J�֬��zhxh�9����Ǥ��J�$Y���t��"|�]}���A����XoI�� QG*m�^'f�;�e��/V��2��у���
^(+I�|ǿ[*�\�	�)�<l"�����x%�*���,���Xߊ^�(����}�L�'o"�M�n��[1!U�����n��*>�eQ�U�o�-C�e�K�t5:Ӵ�3R��n-�.,�+�{X�ݐ����Xh��!i��-mH�G�9�q{#���s�K_���G �+��oQR� y�P<Y�4<<��<d�2��N�ݩ1rS$�wcfg]'<J�޽��q���鷅�s���(AQ���ǰ���q�X��/�ÇoR���UmV�zh�2L�6�iF
�`[��}�f�}"�d	�@w#������}w��&s�u��?E�]�����!�Jg#XU����48�Ю��o]��~m�"C�8���o�>����f��M+�#>~~�����J��n�j6H���#�hP��F����[��|<Mo~ u��;1�Z�����r�㵮�H�C��Q�J�zb�O��4\qr
b̥6���@����[�?�U���ë���[���i��S�����C�D�W�I-��]*�ADS��q-����ܛ���ɱ�3�4
�P�F@y�o��f��i���q��*�痨i���ϟ?�	���rV{�6��b�/�A�\��&����
6�J�[�)�<tOH���t_�n���t!Js��H��;AiD�*ixk�C6!y��ґ��j;�H�A���C�i�WIt�B���h;�+�W�#�#��<�;U%�^پ}�p�������KM���������l�M�gS���/���@jR��뮃tE���rvl9��Ձ�;w�<2���J�Z������} �I8�}���a���Jp�Uapz�y�S
�YgK���]Y;�I���U!�~� $��b�������$~u"��L�(�QM���@*^ �@%�|���VO�E�{q�K�&q�peUU�.1+�eH��ׯ�S[^�A����4a0��Ѷ�3Isss��I�����n�U��L��dû�O�K`
0�[~��Ͻ������Z\����3�J�C��ի߄cy^�a���5hp�v/$�һ���o1����3>~S̽4Kv�kHK��<����u�*��K{A��#U�,q�A��F�p_��/_�<b��)��yqG���l*7��!S9�|�3��M�Syyy��١�6y�Z�l�aY-p�9��(�c�Pu/P���a����o���:>�Y)5��+�����Ӭwi����{Q��7'v��:+
�`��e��I����h;���q���bR���ה8��h�8��Zx�2#;�@{VR�|L�TJ���ϰ��;�`����/�,(ƓwNӅe���.�������zw'��F�@�]����&�п�E��K��bYk�m�=o$~�v����Z���|	̙_4(l��]P�gzf(�5O��]sp�<A��_+޿`y��mb[�Ļ@�H������1?�Y��xC�T�8I�{����j���V|jii��"p�Am-����`�73�e�M�5Gr�k��)װC�(q�AZ(���IF��X?�����ڦ���ߛ�znF��|�T�jm)/݅(��oPRk�ǹR�)��-�.�m.�N[��0
����3�}�3��SS�S���sR������������Ġ��x...�q|暰|�m���b��� i�@�ZE�$��T\�}m&�յ~`�/��؎��[K��HB�����6I)O����[a� �fW�9X֥��?�K-�0��(voKB�C�fa�R�¢"�Q����X4-��/�AFs&d������Oi,N�����q0vA�[S�A7@��������p����T�Յ�'>��<�%����	�5G����@�^��簠�Ck��R�ხ{qϩ/�&��ri��A��A����o��Z��A�����e���t��U�Ty7}]"�d���%E�S$�%�� ��ڦ2{ %pC��y��d�ɓt��x�q .��L0�sw���>�I��ܥ!��2���s_�{����Z���!y
��c��d��v�TO!�(#�?~���q�ѭI�[�6�L�ي��x�[�2���fп�)�y��(|*ۼohx8�A�{k��B�H�3 ���ݢ��^>mJ-���n*�O�����!	u �&�8�ꪑQ�nkF3�Oy��bV��|���w)��]!$^W��_�ے�x�Sm�����ʈw:h[�q��-�d���4�c�ǌ+��XI>v6 s�>	��S�!��,?��B��'� 'ȴ�@W�3����?¨W�"ˎ-a3�6^��i/��+M��O ߟ�,��^��A`�&@{�d���]/��*$�����z$D<*y��Y�]ւӭH(qy#�)8'M�`&s�,��s8����ȐY�?텽�cz�@�T�'�PO?�N���da肝��Ŵ����SS]t�L���,�_u�ЏԳ����e������rM��f�!"����L�~dd�{��ٱ�լ�N- �gK�Ր�$v?|���ݔߤJmVUn�9���T�j٘	�7�n���c��~�[x=�����P���0{�g\�niS{$<�e��|Vv0~L�����Q���]^ᯥ��:�Ra�T��5��2x�"n���9�LU�cuʦ�eQR��(��?�J]ȗ8B��Q��]mZe�nVQ�F��ֺNj7�c�!��,$�4��H��ߕ�0òw�2{&�)	Ԏ�`��T�J7D��������A���(���G��HH��f�ڙ�/*DxvԘ� 7G���B`�w�^ñ#��ުQ�QȞ1S�=Ȇ��.������t�t����|���)��2��݈� ��8�8oEi!ߞ�q~c��g����:�EJl�}���~I
w{���٬����F5�E�T���ʐ:8dԬW*�c�j���j{�3��'��M�j`�cY!e`��|��L����y��ל���Z��U���VnOCc�:��p~����4hֳV�@��{��Mf��& :��h�Ε��B║a������O#x<��O�w���TZ�������p(yf�l�P�X϶��`���A�3U�I ��:NX;���W�k���f�̓��Ntip��(�/��<���S-(�
��>`�N����R\xo��US�T_���d����FPd<�-��zA������e�Dv�O�N>�/���iS����O?�aV[
�Oŗ��DY��Y�_6�1���O�<�E��ւ��ؠ2�[���4ogI�ߖW3Q4U�O�;�-�����b�t��Hp��r��Q3RQ�3
�]9虙�%Z��*p��3�B��S�
��@����!aaR�q�0K�&_��f�׳}��|!V�K��M���1�K��!�HR�VL�f��̯�(&�ίS�eJG����JFNJ�R'=x\U��M<n$�9��ms��N��N<ם��S$�Rh-aI��xb[���:�+�� �za�����ê��*���i�ղ�x-f��w��t��MX�$�`�L�Թ*?�(wJ�,R���s;$�e�qr������
Y�^�s��Y����G�=�]"���2e�]�j��������z��.��@��p�l&��SC����q�
M���V�g��I��� �^�E��jF����#[aV�*Z^�l��8��v&}�I��	�� Z&p�f��L�\��̖��7m�h^O5Ͱ�Ɨ���M�Sq�G���Ŭ� y:4�ߘ���En7�������FIkf�l�<������\�;�Bv]��[������G7|^���J`g�.	K�ӟD��8q�x���T�-��w+:��-+K̊��D �J�J�|��0�@ufP�,�?ڈO(\�,��Zȧ�c�gT��ʖ��^��[w�a�K�{dvB��u��E�Y�O�X��\Di�:�n:w�ɗ��ʞ���֖����O��H�/���
�|y�b?��J�hp��Hh�@?����,��>ګJrQ5�7;H�w����9.'S��hs��1g�"T(�q/�Ka#�e�I�֬@��@� �ݫ���n2ȇ&A%��v��]��f~�i-ٞ?�d����x˱)����G�����D�9T�i2U��l��9�Ւ��^ \3m�4�'�7=�2��\�R^���6Z�,o�*9P���1���Hq���y�^�d3_D�'Ee�kQ��㚜�.���:��v��8�M����Vh�B��R�M)���;�U�W���u�9���]�l�=g�IɎXD/�Ӽ[Xi�"�DX����5G�\�!s��K��:@�$�fޢ�Σv`��y�!rӋl�{c��o�t�c2+1m[ޑ 'I�U-�k��6���wM����iR1�гFUI�MXC��5P��N3Q �}>/U���X4K��K��	�h��&�� ��v뢀ڲ��@�]�Y8��0)��-f�Z�V�����E#i��&g�{_�]Y��Rq�z�{l"����!�d����ʈ�~c	�i���oIO��`e�Yy2�ɪ�n7n����̳_�
?O�T��5(7��?�2��X��E�ٌ�a��]���93� oS��(���ń!)�̞��u���Cm���%V
:v���&=��%7����'y `f�1�z[j��e�}FscЛ��M}�����V\��Դ������d���˚&%f�ӑ���a䲎H��b��w.�̯�F�$�q�$�yϔuQ��b(4��C��dU"��
�b��R�����sr�q��V��7��?W'���s�ϟ�'Q��Bc�bckU��fkkCV��u��wx��XA`:���Q5����gEbM)?�"�&]¼��]]��PVmE_��i&Eh�n�"a[V���'%�/zU	yD���I�CIn�\YG����Ls	�49{Gc{h�E��2��(��n����x�����!�5���.��s{/��n���p"cϪ��͐~����C��
B���<?��~�kW�x���ny=\+�r�(zxM}s�CP:�ϛ�������KK��2��b!�O9ҏ�p-�AξQ͹��|t���j�<�tF�q ?�.q����a-�sJT������kB�͟g�}��K��A��[�3���J�
H5,����M�=J��4�$N\��L����rT�w������zj��2�)�r�/u���eg7�u�1��ng��\7�`U	'|+%[#�
aD�]W�,#���K C�;09�~k^�����>Lc��H�n���ޙj�������Q��1�EV��7	y�Hl��x�W�i$�}x��՚�$����TeÊ/��M�!K�n�:ơ���"�
���Jm��#�1�~�p�@�b��cR�X�X8��._ҡ|։Y&�% ��|k������lǄ{��};Zm���疨��YV���x%`ɘ�f��BI˞r�,��/Jξ̤TӆX���e��q"T���B��u���[��o���D���Es���~V��k�ۦ@��>���Di�����	G��bl\���j�J�[픙�
�04�I�k���~��hX���x�|�i�ϒ�V	U��Ɂ`B0Y��X���Q��h���	%3��5�w�>57E9����j��B��S�cs��0T\t�P����˪|{=D�3�LҖ��c�0vZ{�߽!>i�8QLX��s�S[0�VH�����z���?knn�E��ץ�9�;��$�o�c�I����9�5��G��xצ3yx�z��������#y�Ǿ�y�n����kQr0+\������,���=�@9�z����_��r�l�6W��2?�ӻ0	W��ߪ�3}�***��y�w`|x���Ws�������hj�æo���\�:�����A!�SLm��;,BcmF�.]��!�/p>�dԚ?�#M��S��'�T���a��(O�g%{�'�S����U^���q蹅P9TsS53����ؒ���=b+�0�n�#T�$�*U�Q����Ȯv�n��ǜ)��Kh��r���P�����ٷ,��U�4n0Q,�	"=�_����&�������Z�U�a�3���-��_�og���3! �ǻQ���x���*w�?m+��=��v��҄�R�_d���Z'�2��q��T��m0ٝ�OJ�|���\�퓇"�4!�V@�-~���8ʅ*K��v�m�:�fl�7����6�PZ��|:2
G�I�.��Jrݚ�#Z�#��H��a������i�q�N-��z��e�$X�)�r_K�W�@�"�dz੎�����?�O�>W%�n��+�WL��=��q����%���Zʻ�BY��M?��ϙ�ϯ�O��m���t`J���p4��a�*�7ә�#�ݞ�<��1>�F�ULY�<�(+�� W.G��4��񚩓i�����=L�Z��287E'�Fhow/M�صkׇ=>`z4H�
A�/k�����X��i��#��b&#�,�Ͼ��-S�������~V���}6P�U�4(�w�ﺥz��֐sZs��֗��]!�%� �rrru��+P��	To[A�����\Z=�[A�D	�b�uW���(�6�O��md֋x����lմ��a�g�� $dp!r`wS$_����P*ݔ=.��?���y�w��w=�8��O
�ɩf�w�9����|��#Z#�Iw�k����m���J�I�-D�>(9M����Ip�S^��T�irz<�A�g�� <���_eJ�ٿi+�B`2��?��{����EgQR�l(�?��I_{�#VI�Xu4?P�奙	U��,���
��x,�d�<b���K�ӡ��D���1��;|ϻ�E�|����J������N��>smF�=-P�iKjvl�ó�>���G��4�q�̏S������ts2j��{Ks��N߉μ���~��
ٚ0�7"���+��o~�΋����^^���:��=��p��pyQ����^�ޢ��,�e��0Gi�]���N��� �_��M��&LG�D�;�4�`^�P�Y������h�[8���$��tx�2���YB���ԍ��f��U��<`�xt1��$ߣ?<i?�)�Xtn.~�7^c*�;N�Ñ)��Ս#�@P5~�6�X~���h�h�3b[��i����!RH�ZPB�{����lu��T�l�^C���R��9��+s��o��hYA�`�`��
:��}5��5G���C^7��J~�ی�(�ݞ^�>Ѕ%Ш���\q_/���`
9�. ��&�Wρr+Lq��o�މCS�Ķo��j�x��*#���a˥_�M��¤���/�fef!=�C��/sI��s�G{���s�s��{#���[a]?J�.��$l�a=�o��_����afg;����P>�4�1��g�Q	�]�ʳ�����F�{�8��`gg��Oȉ�,\0���Rv���wg����K�j�!D����-α��2Q��vg'!�������g�|�Iw�]w�[����7�|v��>c���\�f������h��Oފ�Ut���gNK[%(?y}ՙ�(�9aWCs�>h4-[J{�Sm�U�}N��f\{����p����	���a��L@h��j�uT��-'�W��,�y$��*���_��.S���x�lykq���d�b�X�4�V�?�'DF���|xA���c���H{�� �:�kb�"���{�[y^��;	��zXݬ�h_H�f����?�(�+vظ?��ך���Dn|��m���b��JRrE����4���S�������A�|�Ҭ��#2����T������*+�E۫f&^��
B�XVr�m\�L�*ѿ ay6%���K�bUg{�Vqn�^��QVfT�Zs&��9z�[gU�����é��c���S�J����
jw�uJ=�-Sfjt�}��~"�M�w�0�S�r��X�r�t���U����\5]�aJ��){TY��oN�n".`�+4p7e]��!$�����0���3��$���}bm��EϪtU`vF�.Wn���9ӎV��`�;{�﯅�?P��
��^]��4x��T#�>�L�U�c]��o�w&	�G*z�A�I�B�����bWt�XO8��9�,?��*WMU�Ȓ��'߾F�z�{U�N�����A����s��۸ڹW�Y@��jy��*m���d��������YXC�d�v�Bs�r7B���:b@���}��I"��?-���Mޟz��,���ݱc[q!��󷽃��A��&K�:~�^y��0��zT��cx�&�<a�i%�+qc�.�m�-e��|<	b֕�@yDAg�
X�_~OqM��p�t�N��c?���_�����!�eW����̯_�[���lpX��n��Y� +�z7E؝U�*�V�ʷk�Lh�7��:�E�&���"x+�&b��T%U�Rbx-��Br�?�p_���K��,$�|@���1�0F�=�Χlا�y�/��Q�g��5���d*�~���O�J:�ޥ�ث��S���ga���4�#���� �J�]�*	�����gj�1e~�;���e�����P-�������NE���ϟ�"8q�Z���
q��##���F�C�y��T�8��"D���Kw�����ذ��b{��O۷9|[8s,u�[۔	�P�Vib����Z;�;?um;��B!A���=#Y�*7�0c�E�2���{��d&�&գ����Y٭l��F�<C4Ԃ�!�gt9�׻|@���K�{�|�>nZ���FZ�ު�<��M����S������HN|���S:ZZ�����J��D�m�������X��%��Zh�(-��[� �$�,L��q��a�Eno�'M�A����r%�/_�Pa�����X��,���14�z�L��_	3�
GBc�9�}�2���S���؉y䠗��/0P'��YS�y�@�΋��W�����b��qc0�*>
R�3n��S�W���%?�{�o��	�p`��|dlaa��V�Ԭ�)E��t��_]��P(-hڊr��S��7.��i^�*9�:%�2��N�"nmSn�58躻����ܺ����.&�-�Țz@�e�^Nl�=vâuv6ׄ�S���	����n�;��ϲ��I�����3����O,~�r�"�#�ڮ��N`��}�I����8�*<u�L���U7�S^�j-���9a�2�A�����si�Ж�T%�jֵW��
��������֛lWf��9�T#����%�$���za��)֊OG�\�h끌n�>�r4M���W�׻5�c�l��u[���w>�}-����=(GX¤O�������W��ڜ������<�S��ڌ|���Z�����#�B#o�e������v�k��7S��|]XȂ�%�,R2H��r�@��^[���l�� T�����n���b��U�y�7����O�q�
�׷�+q��aD�w��^��C�w-�	��9�X��§4�����s6L�&v����[Aj�u0�w�eV	��ʆ�.��X0d8/FV��,�<��L��E�.w}�ڜ,f�k�!fM1�_�܃�2��Ҋ�fQ��t�5��d�ن�s2��.T�5M
4�m� �6�RP��Ջ{��llR����ŗ>n��� ��;���f���-�1��K������|�y1�(�����z�31�S���1b}��|�@�����V`���ֺ��`�KG�o�@(�X�F�I�U�Y�)F��F<��`BX�j.Xq��>�B��f��=�<��Ԋ�_@����i�L�uK��6���p�]ߝs��՛��7�x��i�!'�RjJx��%����Zg�2&��.g������VffZ���}lBB��_oaw�4�^xg�Tb��Eh�I���E�Ů&���cZ���C�i��\��+R��+��p�����h�����i�}�J�Z��C~a�D�����R�N��A�����Χ4�=,,,:������]^���1e����D�v�ι����=�α���%�����`;�=��V��5C�V�m�oo�Wi��ko�f%CW� `�P�B�r(���I�o�a�ݿ>g�"0|�s��d��Fd[W���V.m/�]�wh4Rt��R�����A��ެ�r��l�߯�U3-a	�'�B����RSS���������}��uQ�^���cc&���ס�4 .�.Y֝w�����(X�!���L�5�����Ֆنd��w]
 ��?��f���,t���R ��}=/+�Ɖ3#��I	����k/����q�Y���Vݜ�5��X�D�RN��|g����|�_�'k���1K�F0�zi)���i�ӻ����J��xv�eO��M���[ <�S���!�M�ϸ�f��)�M�����=+oy�}�$���9#���γ,^�]ap3�1�ݔQ&�t�q�_>�: 6%L%f��<#�c U���\��`#��CkA�lV�x̲8��%7������"�/��mϦ%�հ������}�.���\� 0d3����'?tp�%P�hk�=��7[K�S���,��O�R��RpO�
����� ��˥�|~9X���;;��$�����R9H���z�{@;B�\����<���P�up�O� _�,��v�Sܻ�&��5��LL�fH�n�� \#�)���y#��n�@���gIY�z1��|I_���ye�h�}(ZǾ�w����y˯#D��H#E�A�&�%z�k��''�l�2歐2�	��&���-8ǒ�Jg��Kc�~a�c5
�o1k�7���!����%��?js�*�n�����I/[āMD#��۷?]y��~Lk�D��q7Z�R��$q�׷Ma�@pM@��U�����!���xJ�~���,��;j���:�����PM��MS8k� ����ۅV��Y��x8qm��E*FN� �(d� p�h��vG4�P���J��S�Rq���yUx���UV��Y0�r�`�~�5>h�\L� �~��� �1��5H�A���h��J�P[��\����L�B��3�+4ӱg�o�+���d\hKt`I���~q�z�u55�e��-��8�J �����:V"���?ȍA&��2�v��i/6��Mh�E�pU ��_9��do�i�Un<�n��	��؈� n��*����V�L<�B�G���NǗ�=��[��v��Պ�!;���p�:�Pٟ�P(x�l��K�7<�����i�
0���:�֞�}�{���h�7G_�l�Hg��?�dE��Ç��6o;��qs�k%�Uj��Jom}~�-�]ɱ��69%ki���º��Ɵ�.z1�(�_Uç���>�F�Z�W�#��T�G�UXqa�Ǩ�����͠�r=�8FxT"YZZ
�n������?&������Y=�A��	9��던��:�ʬ��/ �:�q߰�5;ui��g���5w�����&��UI���w|�"�n�&u?|��,���)++KV��5��v��g�{+�(��a��[�M��r����I�_���CP����M��|��"�3UC!�$v�^i�5��7.v�(�SI�c<�����$���rb�A��w7Re5`hi�`|1��O��V^�pl\��Õs)�n@R���:��<��B�QD�̪K�?mt�G�k�oq���65��C�vJ6p���+�x :;8+[mr��C�3P$<B�_	��r�MD�Jha39a/C �[�b���
敞�$�*@�v�nn��bC�}�������s����8�Ř���<Z��q�R�]݃�� E��脘A��d1æ�G������8�W�U9В��vv(���Q�@RI/d�w����>m���Mp�$��֦0�_e�1�Yx�jk)=r�ު���[�J#�Bk��ur?�Ņ�Y=IT�'�`C7�s�]||U���[u�hk�T��ֆ�g�c"���Zn"���[�0`j�/2Z+_��uE8�fx�&+@H��d'��u��M�y�����8#�z�N��SM���'�L��E���0_ ��Q�3I;���Ҟ]�ګ���,���U�χ�T�V��ŋ9V7�s�W-4���w>��	���L�Nq���-�1*�k��614x�B@*z�hY�`;�j �砉�4� �Y4��U"����NtHKéu�o��i"�?v0RCr1��)q�{�ެѱ�b��.���2%U�3�0�#��f����5M.���S� �v�}�.Ũ_��_�E���B���� �W�h,͛U#;t�xW�> '���nD���V.���jj���_�EQJ>|���ʜ�
(��|\v��2H�'�2�PV�0&�f`KO3��s�K綗����A^����_CϦ�N>�Ry��>-[m��nݚ2��Qz�	��/��E|",��:T�	���}(�|q�$}��f��U����aЁ�<��	��gϞ�F���1��,d{� P�ak����B�`/�8�"��o��������:V�� h�d<Њ~���8�zl�"�ZLh0�e�Mo����{ȈW EDGE-����������>}�F��J��E0[�ѐ��w�tGH���)[K�i=��p;
J�~6���#A<Zɱ!��~��6��Br�fC����G��<Zꘓ��@�?�͐)#F�7g����S�r��� Lʒ2�r2P�	I8n�����N5�E�O�%
���D(�=#sm��%h��O���ww>!�9�Jg�h<�9�YU��Q����-����m�>pW���,M�bt2)�����T�AVV$��I"���H��y�� �����~'�NWd~\B-����A
c�.p��onbԤJ`˯�6��ʮT��`�ʊ����nm�׽ks;r�Uc�wQȝ��eQ�R�^� �a��@mZ�Ǐ22 ���f�4%�����9���s.Dg,�IjW=�498B��|gy��/gv����}�%$iuׄĻw�@Ƽc���O��#�v�*¹w|�)���O8�|�2**���^���� ��9L2	����s�'ԗb�[������L ��t���m�Ɋ[�;~S��E�h���!�}�����JY�Pk�z�/����Y[D)g8��t�0jJ���a���B�<��#9�]�~�2���q��G��U�gQN��~���I
P����V�s��=�h�b`��Z-�*��'�)�0p暫��;1��P���gc&w�����k�������p��Y9<�g��ۆ�i$ZOo%�� ٩:))	�a��(���;�Èn6~��C_m����Nw��Y��8�����!�&��]�G$$d��F>�cM�pd{��^F�W����5�zԞ�cd�>̞Ԁ�y1�e���P���Ǐ�N�ǭ՜@�3@�R(���|5r�W\96�����>��;g@�����b���z��.Z�����!�J#hR���^:1i��ō����kA$g׫H��YD6�
��p�D��=*�ZD^��N'�0�ݲ[�`�_�Ɂ����6o%wtt@ (j{�����KX�{ 1�f�V&_�hG���ȩ�m�]�~�c�0[�Mr���������Z��r��i���_��vHLc���/|!z�1��+�1!R�S�1�M�
x�`q��<�������h���j��l���uQ@+:�ʛf|Ĺs�V��������[��ϝ@U��:�YP�M�m�������P�pR	����C��*�%?�m���AKG��0N|-�;8wlHj�[8q�mm2��� 	JII�mLUKL�l�al�>6"(ʹ��M���\�`h�Q���-��C@+1̀����.f���)KM���:P;0�e � *}I2����9`��n����xP��Y�\��:r�c���	���.��<9��M�
���0��얕��cW���՝s gmሥ���6���-���� 1���V"�/�mY���_�Í@�&�w<U��ܳ�/���b�3c{"a�7n$��Crઐ����tƞ��'+��1������O�lW�v���q�P54G�CƁz�B�>��1����a�o"�m��,��
�BJ�N�Z��JS���|�T<Dֆ�:�'$<�μ�{7tl�wz\Mۅ�Nw������5cD�J�Jb�62� `�f�ՠ���J�*�2��R��m�f��Ӷ:)�2.��s�	�D�=� �OA�?PO�6ܰE�I	�O�t�f���w<F����e�e=J{�`	��2�geiY=7�V��{��V����SV��y�ӌY�_�|95���5�4���{3��x�N�6���!�#5j{@%ܭ�³!)����5u^��wE�~�+_��������C�9��9}��J�(�z�S�����q���*�j�W���\�#X�;��˿�l}w?4�}� A�nSt>5">{#Ѻz+y,�xr�����,ݏQR�KHDf�C~������n������n�-y���F�&�����ˮ%�����daR��ųsO@�	���\���_�8_4A��0L����!ن����E�����? e�=�{b#�=X������P!���ǰ��,��I�ٿ]��XT�fgg?�T�<��a�ʠ� �.}Y�r�6��R[������CI �z�^=/=�������h��$���߭첲x?�#�ːWz�lT�,���y^v��(���\���SyI��9�ak�-�4W5���G,d@����Es��'�y�ůQ��ړ��@��p�N�&w�~.-�=a��.ʊ�&`&.u�쇈f�+���(�?~��U�Y�t�@;IF�����UǾ�e��I8�L�Hܦӈ����n.55�p���oXƀZ����2�:��܌
p�=W��o���I����𫃱܁	3sm��X���IVsgY��cS�R72g���j0� �O�p�]��ҫ�]XRR�g�iQT0Fc�����Hmmm�3dee�v���+`ԓ���쾬���|O`�"�"��^ۼ�/����LJ�v1o\�����������ԕ�'|� Uo3]�¯�@��ެY�.+˥�E �lލ}w���	�[��}�&��+����/�ۀ������I�=s��K��%f���<op˵k}$��>2��+C��v�c����i�BKY��R����>��	�9����8N�F5��8�?Ź�(6Ѭ�$x ���˱�
�>�XˣtJ?|��7�����J�^)Ֆ �ĉ���G�1������CI54��	q�������������B���o%�8�,T
:�S^@�t|f���8��w(V��Q��D\my �9�R��ح������k�OX����hK5���Β?1j�l�j]&��Kr�0�����v���ZĊQ���'4��8��=t�����2�L�ؼ�ƂN�tڤ5ϫ��o�{,f}�~�LW�Z˩G�:Tol�q�w*��+��tm�ݓ�Qۛ�������Sǜ�n;������|�ϯ�"�|������5) �gP�|�C�F�ǳ�V��Ro	�pDso�L���ZaR��!�ύ��P�/�_0�=�-�'�MY{z�|h�7�
��J[v;o�b=z�n��|`僉I�^�-������$�Z��A+�g��12t:G&�ƿx�@!϶U�v23�:�e��-Ӆn�'�l�l����jR/k�� �G�Yv�uX�w��<L��[�+�j�vT;��Pw׫܀%�Lv�B %X����ɏ6�	�`۱��r�����㡉����Wr�o@NV��~޲��|9��|I�u��Kw��rͅk!؁y�@�;�D�9qO��x�]_О���ej�>��^�f��Ce�Y��uZ�Y�N�z�~ {�1��D�!�m��OT�:�0�-�O}�:��`�*+�](���
�ﾔU{�a|�t���:�w����)g�oD������U(Z�5Q�����Ui��)?��G��k�~� !`;Q���F�K��d&�YAb�Ԗ��ă8Q���_�MD�2�X�}�՗�4`6{�ܤ�{x�A� �x�fkи��K_�fW5��'�_tI�y��i?�p�J�?ҁ=wJܺi�7ϳ�[sz2P,�U	`*a�@���	�8�<�pb�e颃������+�/�й���ZS�G�^�z�vb^�t�_��`߼���eq�ѳ+�/ج6��,�@����p����}���"a>�I5/�X��W���M�;�}��Y�1I���1�Ţ�vp>�7O<�Ϧ��1�ژi0��z���?��G���������c�l�/��G�����S��vڟ�⎯����Q��������9d���D^;�J�������|������<�o�kZ&�������_�/��K7�6B)�A[�/h讠����@�P���}��g�J- �^�B�6~͜�P�X�`9C�i���q3p��'þ�	e&�xb��2�߱37�p�Qt����كI�Џh�?e�j���Mm���ل���I_<�`�3saoV�h�e{�ɼ��]-O-W�����հ�0	ߝeb���vU	_>�]�2��8YL��:Z�G�gD�w'�� �c�o<�G�`a�u�xV���n�cYhe��s��r�:ߕ�|t3�וo:���U�wa���d~o�-���.ly���gWT��z.ݷ���6%��Lɇ|o��°)*3���Gc�iP9װ��#S	�2���V&QJ���Ut��kv`�[�����2ye����
�>q�>frYn3a�7���ٵgΖ$�sjM�)��2�u�늹����bK���yE�Y�-M*��^�*-�����k�/w����G���?_\�j��W�9�+#�k^s�:��K�Ŏ������#�]o��wP�e�����x����H��H�
]��u�k�|���#(�2N3 ��0�������Ҡ�����L��{�x���oܒ�rJ%���J5e��TR)�b�(��3�E%�i�u*E*[�)�mB�uƖ���e�>�g�,Α~�����������i�������z_�}���G���)��d���$10h���|�мM��v��9A!��Q�i���(V�7�^��ϣvYN�<��mڸ	!��s��4�.�	E�\<�dA��^H8�o�%�$P;۾Џ�OP��2L_�Oh.L���DJ{��c-���m)�+��f�)l���\�/k=��&P�P�W_aV��F~��K_�N(��´P�˸7�A����&)Y����6 �(��ͫ ��H�}��
ӹm2,�Y��9��H�}M`E ?TeZ(b��h������J�s)H�������p�b��X:p1�b�S˯\8��w��"	`�&ȸ2�q˧�o��P���Q�7�!�
�jQ�B����J?��B�N���ݤ�ϖ&�����X��/D[��y����:��ꍖ� �,�҇);%��%8`�;�����g�>}I�`�'9����N�ǀT���C�|�%��i2��@2m��3�ˎ S�f���&��G�B�	]I���k���mOd���S��3>�~��b�5���oTo�^8%S-����Ya�ԫ����D(2�~�
`������7���@I�G�Y�6}��`%��V*Ӟ�h>�(�=��P�N1�	_�A�ΐ����g�,L��]`��S��s|򣊸yH�eqA ���S;��~!�a�����29��0k�Zim�Ef���S�4 ��%����%~ZP$�b��T`��~5VZ�o�O|Ԏ��*0hC   ��ڝS̾�`q��hq�{K;���~�wp~�wp�o�'i�_�|�w����������������������������������������������������{��m
���s%�k�~Y���5�?���HCW!E���p�Q^4B6��������uGV~�@Q[<kUf�4G�3��s��6��iD�O~}�B���C�VJ7�H�bx��+P6�Sc#��C9�ъ(̋�Lg�t�h��FЇײ��^�����J�ݏa��\�Ջ�I$K�������TJg8��� ��=]9rY��^��x�@��N6���2Dxh����t�bΡ��v��xy�I�"Ngxe3��z�57�ч���>V��q���_?�41.����M��o�_���DD]V�tȶ���m$R_#c��¿l}bA �Y:���,�k��5���7��S��mo��(���5J��Y�U9�yb�*JR2�͜�,�p�~����س�dϽ�L�`��;HV�)L���SD=L�)u�\z���Ǯ�La_�H��%�ӑ�TZ��|)UPĥ�6w	��wiQ2.w���f|��X���$;��^��p�z�h'�?Xjϴ���D|�	�j�~~m��pL�a>���jė>�{��d��]3� ��|�6ᐇUX�2�9������-ԑD�S.��&c�B�43��GOM��̡w9�y��.P�p_�2)v�~��rťe���1�h����S��_<�߸�B�	��zǇ�rG�́�m�Xť��TN�E��q��D�$��R;��<2������	y���]7���K+m��# ~�5Ц�����%��>��[f�[w]W��~6k�s�O��n:S0_=�����N�2;'�˲�\���a�5��Hx|6��3��;+OmN�B�s yu>X�.1'j�]^|�ΰޯ,��8�����4�<�s�c�nw��(�ۺ�t� ���H���>-�4�L�sZ�I^������m�u�v��y�4���үc��^��x�na7g�sr8��T�w���������#5U:#vS�q�v��fAL���J�	� ���#6HN���m��ə�ϫNڕ�6��<}�mO;�_�����"���W���ե��h�p��٬�i�N0K��Oy�U(^
ao��h���k�|���T��ې-Kt���r����u���M��iYa���Æ�v�����X�Y����jrS�W��7̦��<

_���_�s��D�Y͆w ͜Μ���K�&S�!��۸L�{�i�����L�a��]���;V���	sl�=��4�u�9��Qng��2�����6�X�ι6�~
9Z?��j�ŚAt*�����6"���J��0XQ�c��'����������"���c�]gƻHb��ױo5O���o�5h�I�OIh�0*�����ϡ-<�~��	��2�o7t�$�nz��P�����EȊ��Lu����S#=�a{�j����L.1x%�J�����cǸ�z�j��>���1n���>p�&�UGU�~)�s���ʄ�u�Hq��M�@8����w��7uk1Z[ʵ��818 FY彌2��s�������j.�"u[[ͦA�%.�+�G@�;�+^���)������"O��рI��3\x=,��~5u��t�*DW�ϑ�=/��t�(�]����E׳��CJ�'�׃�c}L��ȿ"��3��ׇ����<�ZVH�ͪv_HvjŎ�*����I��Tck�}�� R��H��"7�qe`��x��S-�?�$:�a�Y������橫_�X�1ӶZ�g�OA�� ���9=�b}�Ž����ӿ��8~3`L�>�[A�0��e,���렞n���4�|C`��7.c�����4gNU.����b�V@5���%��?8�!S��$�@�D����~�Z��������^[P�$���Ϗ�o�w�G�ȫ�7�\~lԥ����/3�"|E�(�����K��@=� �׆�u�����=3�3'(��BE��)�d�m�S 6$�Ћ�M)# ����v�G�	_���:3��<_	q1k�_��8��P���#���S0���z��:J�j#�P�f�]$��r�ـ���ˡܠRfTZ'�_Dz�'v_��?�+���o�o̎��9�<*�˰/�B�uʸ���t:�H�V�i�FZR~p.hi��k�d�9�[����e�EA�ňA�p*\s���ݰ5�|�V5�J��K�|�8����"��#��B�Ǜ���a�4BsGoP�����"��_J�vm�@���N^-ř������<<T��}|�*˂^�@�9���vA>��ee�r�ELtF�fN|���Q& ��:��,�ǿ�DA~S ���Q�+��iw�ŉ���9�s}Į9%	s��]<l���� �B�E��/��$��*�q�-�9��a�� �ĥ��?T�@Wd&�����-�z!����X�chҙڄz�E�5@Ĥ�}p��ȋR����@
w�b�`웒�j�e�17�S��4��p��wegHF-f����*�@��o 5��@���`�*�o˻~x�n��5d�]�/d�.���i�X��ߣ���"
���jIWM;��K�O\ ���k*�T�K�sj:�p�,�%1v0R!�\�h��c�%��!�-�(mW�o��?A_SHṞ]���)�٥�/:>G�RP����rۆ6��=:|���x�U뵽h�jʫ��d��R4��ޗ�r��w�d4����Rr�;�zqQ�h���ה���T���Y5V��g&�=���qB�)��)|�i�j��8�Z�У���I�j �G�k/��v��ig6H��`�"3J��<��s�z݂��K���Ik�Z�I-=��,����]�!�����íq���`Y��F��Y�z}�ǽ���m�8O�gX�y�k���wf٠�=�II�,?�3
X\��˹�����H��$;tȰR^�vט�7!bbF�m=����囲�x@=o�	b#f�s�/+/ۖ����YC���E�w@�-"�*D��IǍ�і�>����6���qc7���Y���}�	�m��9���)���(D�5T��ܿ��6(�sT.�yB���ΩjY��~���#ƙ��Wp_5Yb��O��x�bL�������m�v7y)�; -�E���t��=��bEE{hi�
�]hDl�c%@��
D��1p��>����;cđ�M}��H}��'OL��~���AtGp���. ��w��{�\���)��(�b�����X���t<�������4��uF���%{�M�4�4}���>�M�:I +my��L�w_]g���f(,���ݏ�KNNb4�B��zg�a	���[�KS�/�)�
,����h��o�S�����������:w�Z�Y�ET3�n�YKl@!ˇ9��/)Z�gݺ9��\���E[�����:���"B81��AS�H�CN�vD��V��gsKqN�Rȋýge�:2��N�_����9�H�*4����Zc��$���$�69[�^h��÷a(�>�dN����O�!��"�g�a�+n�,Zn$�e_Vۦ^�v�A'�o��i��_�[z]�Tq�|�O����.U�~��z���e"��-w�}E�q*�'�J�_��2Rl�ðq�B��GU�sΒ|�$���
�a�(���iU����e���A�,�L��/<��c��ayJ"��J��/3Н�i�3T��]��8ǘ1LF��]�w��3'�H����PA�@"�ɬ���51�'֥TX:v%Kq=��ڵ-�B���$;l��&U1&�2�qx�������M���"=.���p*.]�	�bw
�$�jċڧ���<%7UqtB�;��»�@�R�츽-;KQ5T�hw1��VIy�8�-�c(F��_��2H:�Ŧ¸��dp�l�$�7"�I�W���/�d�-���^wc	(���ަ�1�n-A�^���A���o��f��!9omKC0�ӆ/�a���.F3UC���\�U���i�)ͧf�U�\�iZ����I�g�p�]��Lݼ;.����ʣ�T1�������	����4�� ��!���z�9�%�5��0/$�R*Y#-�e�����F4�BP}s��~�?5jԾ��5Y�U��M�LuOdl�&�a�*��x��O���T�:m[��j�~�J�e(=K��g�i�\P���h��z��g�d&�s�&U��hH޽E���?yaQ��P���[q�-��� (ǜ�?�������n��XzME�{u�J�ؠI9��1	�����D��>���Ɏ��NB�N-�0c��x���ƒc6�*���| ���j� w������n-P6�G���
ɣ�O��8�ml�a@i��Q����ī���^B/�)�9YG[Ǹ�;Y2��m^�ɦ�'Ҫ݃�N@ �TV�l'�'"2C��uM�Y :�m�<����3���sQӂ�r�C�<�q1�`o���0l�5��{�k�VFJ��b(�5�����[�yy��< \)�v/��'�pLǆkiDnҙ���ܳ��(j� U�ޒݓ��&��jS�q�T0�<&��nq{��΋�Ĕ��W�B���e�L/F}���,	2�Xk��v���������L�9Uw"��Δ��n�J���.g��b}�|H@X�B�Nُ&����(�u���-���;�hB��iZ�9������⥖l�/`�GU������v�����e!s��*��H�H��/Fsr����T'EF0 �*�j�;���Q^qO��ф
��ײ�"6���{�K�§���������WxA�"je ,O��Ս8q����|N3�I|1�s��l�o�2�|���v����;Ыb+];�n���;��®�;�
tl���9����{u�j{s��\�397�004�p���:#r-+6{/�ŌL]V��!�^_��Q��m~���:\�2jpR�{��Qo��L[�i; ���u�@�0�g��=�.hF�?ba����P��CuQ�.J�������g�%H�yM�@��:ř��o�/!md�p8)Q�������*3�/%��yۤh!�s�y%�/���y;sNB�㬉�<`�W���-%����� �y��F�+���z�G����@�Yo"i	�.�����
Ԕ��S$�<����/";.�rކo���ګ�{j�X�Y�1)�J���g���(��+�洭�u�'b�:L#��X������Q|��h)ë�9��Ԫ��2/,K�;Կ-H��/���%px�J����w�5��:K��'W��&��X���N��g�	������N�����):)�褫d�F ��<ɸ���`�AKE&��:ܗNNm	o��}����������.���k���r�W�R��������p�A����$�p�.��\f�Z�r��|D�w�(��'����4Ru.#5�;ʤ�Y�O�|Ǌ�:n��z+��ͅ��#��]�;G�]���Q<�qɺ3㷘��a�쥕�=łt�2����?�mݝ�	y�QZ�oa�7��7!=SB�{Y�6�]��1�N��h��ӂ���dj�s�2�,F|f��ݐq��:.�~/��z�����VP�ʹ�:#�M�_�Iu�D3�4�����3�(��:D�n��f�n��)f��!��e
�����Qǯ�-���`���8jf�50����d��t�I8�b����(����ʥ9�P�)mݮ���o9��:25�P��xT����Lk�7�nÕ��`P����'�.MOs�
y���0���P���R_H1�HD������w��^�Bby�=C�����"偒���"Zշ-�����Hsu��I�@I�/$~�PV��sؠ��m ;�B�~N�W�s/^�I�����c܊���ͥT�%E�{�ݓ�	K������.m$����+�D�%ԝ�7p�(�����e*TAG�%T�B�,Q��K��ė*��>��R=��Mä�z��p}�Uw���pk��6oi!o6���t0*|�0����72�v˻P�豑��qd
)���:w�A6�Ie8
�	��d��W�?j�&DC��=���S�D	��(6��X�����̱D�,t^IM�@�&�sq�4m]vn�$q���3��>-����%��0ﺕ(<94X
Cqؚ�*^[4�1B��?_���(�,���{��Hɮ!�`�)N [�}:�o9(�~�丨�f���j���;l\sN��Ŝ�'wʍd]�utRG��W�@e�&jw��� �o�Ȓ�p�\E(��C$���X0�%���k�.(\-�°#�d�Z��W�D��L%���|p�rH�V�׺@z�9��IC=��q��R�9ւ'�w�gC� ˢ��kϱ#4��Ӏw���R	9 ���AsK��8��~��p"��^�r~��&�G�����J*�y����c�biِ�.��6.zՀl�9���L}S��zGvG��f���㨨Y=���)�=8P;Tҳi��������f��Hk�R�#<��.��8�~;+�ь{�XdC��E�bV�I��2���=���^~�E��[`�q�.�G{��Nr�>Ms7a�6�Y�=���4Ur�f�Qn<�h>��`�!������!#�92��VI�>��u�*'�_/D��m�����A`�f
����5a���힡4cƫ�0e��;-�y��{?�B�8�҉���x2��.@�\{�������~�g������>w���\�k�9\F~�E'B�:6����T�_&d*�sZ�p�t��C
����M��!?))�;���}M��	���/�Mw����ٗwiѼ��[�1Ka�6�C����{7��ן�ߧ����>ZIH[jp|�x����p�E����ҳ,�C0wh���'�c{>}Ȼ���������m����"�sE��&��R�q@�8� �gԖ]b��+����U�x�mu��K[G	0���1�A
G��"�dA)>м^��&��Rb��(�ҭ�#l�Ad8qe�j���c����='�%�h>
�y�J�5��@�f#��̡��/m��WΏ5��ug�.�o�UC��Bԉp������Yz�Y��c�/JU�����r�u�Z�����>���x7���X��ŏ��qW��P��3��E#�4���0^g8Ҏ��Ҽct��Ls�E�)�h,��j���ewe�'>�=���?���w%�*�C�'�x%ځ{�ۛ�b̧?�b��X�DV(,����<S��zW�i�46�0�M\��o��D�>�e��33�����o�y��e2�f�W�����R���q�鐎!���M�^e:wWV,�l}{�w&������գc�{�aJ�{���VH� �)0�繯�`O��_4zNZI�?N'иi ��� Z�����!>�ɰ���:L�M������ûs�x���2�����<�1��"?�C_+�"�2\���Ow�-ǹ�0��̡���0E�V[@��ǘ��ߓ5�)�|!��У���&YT�@�X�%�-��-��d/o�*lx϶p@k�l*�e��/o �Xo���B|0w&>X�Ğ��y�b�0�#	X�����v���G�NM k�i@Й�QI֘�X�O����
��4�Qݍ�\����S�x%~"2 �C��U/�<b�Rǥ-�/�7����_%{ջjX~��3'މ��*>���/���%��mg���k'|3�k��d��(qs�H��T��縨d�e��&���T S*�����6E����j�/�� ]���������?��N-���Ŏ����-&n@�U.)4ShI�w���Q�D�+O@��
���6lQk�;y?�r�QCn�ܾ�*�����ȶE*��=�߹d�t�m������$�Ћ�G��+��x��(M��8���]�Ǯ�)E����Q�Gح��#@��_2����yY�}�RL�7x��,��q��I�yH^_z�iA�eJ�e��L���D�������>��oK^�X�Y�"\x�I�5�glEwe�ͅ��)B�]U3g�%�B:s#���|���e %,����vձ�p;�0 �T�y��@EU?������3)v��V��4�C�V�@�L�	��7�I~����奬އV��ND���fe�$
��Id��M6��[v{�2]�eH=����e�L�:a"�e��qQ)p�7
卫�>����/1��1V�Ά�Z���)�ÿ?N���k�ȶ�.$S���+�i�=|�rʜ�N��ܑ�X���f��%�O�'�y���D��e�
�c�2A�E�Ih���Rs��lM�"�����RsE�!*`Lվُ"+�����c"���aA2��==�q/����U��2n�\�{U��9?�q;�����V��������ʊ���9w�_v������ʒ�~
���{�oi�?�F�z88�E҆�	� ��q�4n�36�q�h�`�10�.?��L+����~/7M����@DD��A�����Cs�KY/����2u��@��V��'����8��J����l��"=��h,��JG��#�hȂ��/�ؖAM4�a�#�#��j�(��D9RM ��1I��$�.���1�Q?M؟^$�����o"#p~���p����u��!i$K�X�O!�RX*�=�'.�)�R��#��;84�L��`�۷x��^XaSH�Ta���DT7٭Ӧ� ItD[�~�fagط�����K+5P�e��R�-�=a<���Q�D�$��	��
kl��v?y�����y�SZ�ea�;���-�ha�v��.�x����G�#�-�4�`��y��J�n0�o�H�Ⱥ+jD���[��5��(����cc�A={A���:���HKD<N8�IͿ�,�c
�L��|!;9�����C2_i3k׵u�L�B�ք�NIe]۝�2�KYk�K!�+���7��^߆b'Y����tCfdA�!9����� C��=�	i����joGp{n���<�#��솣(Z��w�a|:`���k�~�5���%���j�Q�hn�b�mD���d����DF�f�bD���>�>����`��6�2�>��!) �Aݏ�����~J�zV37>0�4�DnyOV��<�6q0��观^l=�3��v�Md�����(�f��D��<^��pi9��Lj�w�	O_��?�}��y-�^%p�ڋT���H�G�������}�q��a7���`�NH���_��
f M��Հ&|����b�p����+}6���]Z�m�,3t�{���9��&�0��ɂ1��D.� �H���`<'�N������U�Xd����s~Ặ�2�C�� egJ/),EI��.�l.4���"9��FH	����Q�=�<�
qY��H�ߩ��<���[ۭ�kW�R�o�I�r���E�������F��k���=�q���t���0��	��7��#�#�f��x`���_
��([M��ss 0�=3����q/�;;Z��~.�� XU�|Ax�?]�G�塹��f�w2�0��ć ���A�(�&h�9�H>�x�>m�JMT1���޸vM�gH�`�J����?���BY<K�ё���ĴIÜ�m��;z���泏}L\��SI�]�Ď��FD�����o?���Ə!H^i��'�^#��=�\�����V���t��V��t���*ZH���*����*e7���e0���˴�r�?z�]��!��D��Mz��V�*��<N�^�4�9Tƥ�O.aR
��*�A�hI� �=,
#� �r������m�h�n����6Hi�����w�7��|��Ț�oonn�<�E�������z�^x��-Ýek{3��޽령Rn)K��(C�Z3��N}�u���q���_ļ���2˅�L*���b�x?�̬��#�1x�z
ű�F���b��g^}ɈZ���Q�{1��Q�ⳮ�9����N؊����Q�	GG������#���%ƿ��~���[��$��p����
�09��l���A�1m�y�o@�Y��������"����;_�-e�KL���1>��ړ� `���Z�v';F������7�����kV�A��9��PdR���`�Am��ɲNN6�Nn�����Ci�L�k�a�=t�Ui����w��=�����T�֖�-lQ %���L���A��|��Kq%r	�g�sr�NB>����K�I�DSɠ'A2��/l�w���v�6�8}�y�Fy4//O�Vw}pp��Gy�k��i	EWG�����`�F۟c_�`V�54p���`8�����8����J�'V	�E�������{��@��`䜩>�=��>�Op�\WEY��qሻ�cV�z��a��~Ŭ�2��"~[p����J]�"����x�dZ�<~��Q�o!��#��f/�,�R�҉DU�,�9*)+k�s��l�p8�>���p<�������:�杔ɗB�L%���/���!-�x-����R	."9��}}?w�NK�Q.\�����䇬���j���\�����
|�E�F����脪f��2�/��W�X����5��.=_F���c� i�=���64��٩/0ht�1�������8Y�w�ߧ����
7��z��}[F�z:�C�Ο9Ӌ\"�]~��-n��,q��fgeg���<��ݚ�X��ny��gч��蟞�=qB/vGttt�c?��0�A8q�SN^�W�}��+�KVVV~o����g��}|����zj09�Y͈L ��T��<)n���׼�u��C�>��yk������uf�`j i|a��tt?��`煍����+++�h D
_���s���G�LM�������*'2MQ�����Q���&D�=��J�9���'�Ffgee�w�V�9X���>��h����4m("藰+J^�|G�L�e�P�'�_����eP�[�U5ǚh�O���W�ÿ�,����u䘋�t���&k�ȃ�� ʖ��j��/~a8~�/V�����?HJ����M3:�|�� �����lL�Dΐ��s�?i����B�����_�ߢR�`a��2�A�v¤�b�U��V]��zig�qI�n��u]
GU���s��j�ɑ���8e��3m��u��*`�Ƕ*}f�ۛ���ɕn:d�|����9��Cr���1Z�ϟ�9��9�&d��2��7W�k�����Nt@�*��Q"���p``�/t����RcS��&��C��`�B2�d����G/.my^P�����`©����쯥�p�Z�
�R�=&zIkruPgO��֦c��H�B�����d��lȉZ+����П5�	E��rY �>��/w&B��
��� Ͻ��a1�l��S�r����	��g��W=KK^�t�DC'�����/_�{�^�Vk�J9��zȌ[�⒙P�D���v��W���x�Ģv2�k����R��;�!% �nX�Ӥ�/��_�τM��M~���mt�T]<^swy$���p�e���>�2h�.�?��j�����._:���L���^��
��bu�;lY~�������*lpM�>����\���+SI.��72{&���r��4U��+l���>�M!��.���w~m�VU�H���HHpb�e�?3�溇�,n<H�Z�����L$+��q��_����Ҳ ^a}o���H}�.�+E�_C�oY
�B���P�BavC��Wk���s���UNٯ��I����_`(�h�i z������7&:��V`w@���do�H�����慨¯�3�x�#�J�v-\��4�M��oi�Ǯ0������t�[ղ����Ė9�*Şw�{%����u����gWݩ{����Y�|BR�b����"�._I������gϞ�6\UVV�績�����[�B���������`a�Zn~�Ⱥ�a1Jf?VՍ$�]�� ����nXM��tｻ�>}b���7�H�0�k��H7i[�� o��7�2�OJ�-M���O"��o6�JO�l���S��B��TH:>KM�e��z˰�"��'0+��g�u�㷡P1`��m����k�[���B|Ѕ4��O�n�"��j� � v�����.@��7e⽓�Zi� �J���jwru΀��=���aȍ?I�\kn^�g�X���g�ee�K�w�hW=Jg菒B�Q��ل����M̉��&��{�_�����{_�*�:��TU�G��:}�g�I�n;�ߴ?W@����n�YC
&~z�a�^��:g�#�[r�/@���q^{k?E�͊�M��|��n'��^�%rU^]ũ(��t���`w�z�����n>�O�5(��@�����5�:��w�#�"5��C����L��la���-j�&3�[ FA��X+U�)�s=�*6��`�%8И��U����7�J�VΨ�}K�L��;��4s`S��@�T��y���j�@κ���yU��8qv��
�S,`��+�)�J���>�t�k�+�9����v!��SRRR���x�ۧm�s��g��6r�k���h�`��[[[S�q���N���S������}O�Be#HZ1ۜ����@ྡྷ��e{;���C��1���/�����G~��|�?�\�����8�c�̳� ���747;�S(Y$8W}\�1򐼱M���Tf�MM�н���?#3�y�4-��ׯ__P��*��s������r(���������@�Bc䪩�*����� o���9��@���5b��.��1I�Z1-Wr��'��-��Ϡ������s���QC�*�Y��UG�&�a�	N����N�y��U�Ï�{��Y<ӒY�?xz��7��S����p�Tt�����@:�k�`7+Jn`�J�a�W7W�c=�U9iͣ9́Y������{�p�C>�7���`�B!����6���X��̮��!�_���I��1���������8�8;k`���a ����m���Z*�GG��b[[�m��������|��w��SO���� �9"�FLG����s*�o�����k���GH�S�sw�x<���&3:��SY��zj���@
R�b��4ȧ�-�[��bT�Y	*����o1t���@X���=UH~�k5G��^��m��� �Z��s��\s��"q�Q
/��݁����;M��bʁ$��;�KG��|����&l)��啕������;��w���c4��nQ�r=�� �a�w����TǴ��A�"fe-��Ao�������oA���<��T|j^��W����D�x�7)��i�Z�2�>i�%?㪾�~���bm2�H'-w���V�(_wj�9���]�ozNk�~���u'\6�-1p)>�K�`b-P�j�P6$=F�=�V�/��}��ԞZ���ϟ�h�S|�~��3�:�����rR�6
8��;rqs�����{gX���G9* hm�����v��BP@Ab���ޱ���f���L!�tf�	��s#�P�x^]4�n�����+gd��g�Z_��v�K�Ә@�k�;��C�ڣ�㴳�3��tO%r6�P���xk���qq"|�1N��|����/���Z)��+ŕ_�Q�Im3bK���\Yed��L6�y�!������|�7�\)�(����nG�L�}XS!�EDFTX��R����)v;gd�_�<�������nzv6e�,�@r{d>�譓g�^] �l��(.��SI`j�����e���4���7>�8O�x�?[W��g�猩�.�h�dw���O9�ŋ�<�ܡu����x^oՌ�^��[,�e�����0#�:)imu�Hў��tB�����8�Wq�JN=:%���x��K3&��r5�6�N�R��:�s�Sp���Q��L\΅����5������wl���w3rG��6(c��W�Ő��Ҡ��*�f��6w��u�b�٠KQs�:t��.m�&�Z.+N���t"�n7��ߏ=���e���L���?���1?KI�~��O /T(���qž���ԻSR��-��7����u�=>��ΈP��G�ֹ ��L����M��S�Ug������G�&�s�,��p�x��^k�@ħe3��9�yy�#��T�4�R@Eg ݞ�ǳ��P���.��i	���$��$dFH~����s�Ң�������O����ƾ��:��0����,ZY�N��ܝ�f�p,v��]Z_�rT���
�~���?̤��F~�٣�H �����2g��bc������5���c�E�g#fL�3��6���PE->�r� �*0��3b��]����J.�����-���<-9��C�ogtg�C!1����+uoQ[̐&#�f·�B�0��j��� %�6��PǈcJS�t�ڇ.��g���U�Ote�/_0[L�YY���ba���λ����U^�_�Z=�w�!P�vB��GϨ�N�=�� h�k����퇀���,$��ܤ$p ������9b�5��k��i�a�ȑ��ܝg<!�;W�X�\P�࠸����K:a�`j���Dd�B�d�G�w@�ƶ	݈��f�����3���Q���Կ�˽��6:��V��@P�O��O�&%<��g��?{�����'�o͍�+u��}���S6e��
����n>EN]&���QŠL�9�I�YaU��75Ey��ϗ�����{�7��2��㓔��%���O��$���Г��	k&f�ӵ���Q��H��;u0�*/[���Zx�5"�J�G�\
��;lr��@����8u R�TR؀Ϛa ���Ѭl#��Ġ+�A�����8�8���1]:�CRb'^;%�$�W=?��mPJ!9MM;\\R"�m��x�tS�Ё���=��;���{Bq���M��!%�1*�n%b끹zyL�k�kr2�?"�����.��d�U���$��`�q��I�+a�w���.{Ѱc~�M���b�?5̧#Q��̾G�oke�C-:�X� 2Uo <�$��$z\�C�����D9C�J���X�AR92{�R����ѡ�9"�7	�H�'�8���T���I,�r�������:w�"���L/��q��s~�� �sv���D//���Ass����5g��JY�AZ���QU�/.yo�Z�w���&o}�.H��W�	��(�`��:j�84��
zh�������~�v���ڒk�kd¸!!R�n�|�����HVeb��6����᤯41���9Z�n��hzbj����ֵ��=�B��˓P�E�~wK2Hv�;K�2�Ν;����Y�L�*hp̺6�!�3��?����w6X	I:::�[.�R�rJ����[U�`�F(G�l�P)��p�v�zn��	�z0d�g[V���>hf���چ�;`����D�}����|�,���?L��y ���	�=� w���P#O��yQl!��Ri4���f3�n0���7�RZ����x׭j�$FVǖ�"���Ƹ.�%L�>@�_j���L�m���޸���<���_�b<�����m�������~�CW���o�o̴�x/ڒ8t�ژ��y�ڿ�YRR��^)���t�͑B2��z~S$d�ſ�IheL<��͗N��;G[|6��Y�8`~�E)Dxccc��`�����W� �aP����<u][s��%7 ��IW�k��t�� ʷˣ+mX�@)�X2����}�G
tX�����B�(@R,!N��7��9
�Sx),��
��
�����G���p\�re�-����ij )���^�w���3%$���� �{m��~∣��_e��Z�ּ��t����_�#u+(3Oz�6���r��M@RC�t��}�3 �k׀��}�o�)%�`7�{�f2�@B|Lb�N����+���d@L��u�J Z�����H8ܭ�}L@}��`y{��]ףj�u�Ha��w�����B�	�j���ڵ�Z�;�c��٦`��O���R.Z��D�E&ޖ�6�:�%��͜��1�_6)�n[�7�A��Q����t���I�.���?�}c�.����%'�^�-U`L�.���2\ ���um�m�][��j���|I<���)����У��v�u�F>�W�){A�{�X	 M���f4	bȹ�����v�'>���؍�� >k6�w>d�H5ǚ���z`̪�LR�[�uSyyy{�x>t6� ��4��tE����[u��х�,uEbm���D���а���.�I�y��iruz\*t���[gee]3<�����fg�X�����Ii�ZqS�P���O<���A䵁]F���lN���dm�V��1�����AT(� �W?���=V�̗���Lr���Y��&�3���~߫�R���]�֐'�i�f_. �L��9�1%k�����WE�)���umdWN|�!wz�C�B<F�f�4��y�ھ�~S�l9L2�J�&���Wa�RT�X+�Q2p�T��q�o<@;f�X��+�cR�C��C��" [ؗ�VF�@�)���.�h��$I�r0�*Ր�#ץ��m�I����]?�#]F���:e�2�>�G�,a������w*.�,�lVY?�yXl��I��A�r���*7��L�%����<�*JJ��:*-�2�5&��jdzU���jO����33����gö�$[i\@@DԪ�����a�zVo2�~C$P'yxhBڥ�|�e�$���g��K�z�g�xi���_ _�3�T����rg�jE�WPaT�N��%$%!G���O���J��贿�"�wK��nH$,j�W4-i�Xʋao7tS�ww����O��_n�\�~��R�=�������[~e:�Z� 
�	u�����?L<f��V�I� ��y�V�ؐl�ȥ�:r�z�J]Ʋ�?�V|h#.X�L�����*cf�@Ĝ5���z@@`��������$a�=�K��O����^d]еY%�,�!Ց��`��?�-���k�cÞ]�H�p��4Q�MM�6W����a5=Ыe���ސl&�lhmݔ��w�%[�p��u�)Ӣ��2V�H�c&�v����u��06p�����um���!���@�&�|�y�bZ���x����s�+�җ��
זoh�{��f����^�аu�n݃@�\p�/��%n�>z4}�n~h[��Ͼ�j��a'[���\�%75�Ng��юYO$�`ۏ�	��$��2�)�F� �����\Ⱥ6o���l�����Z���*Q�zSӪfn^> gt�j��5mh+�t�e��hր�rؗTu!ҳ�VX�ݺ����H�v_�C<(d����-I�z������Pb1�i�wD�w���k{���)
�HLJ�oooO�ص('p�����5������݇$CK�v���܀�`$���SO���zx�f�i��\G��Kg��*�e2���4_]�B�ބ��V �߉�xJr�Xj���1G¡��� �_ޟ6k-e�iw�?0A�1������V�<� X�27�.��,��5���^��i��{�R
�-ҳ�]��}�H\	�E���!�g$�����;R���)��E_�迄5��oJc�ϖ� gJjA6T4e�����wU��n�Og��ʾ��8
H.�k�%�Tx���������{i�_}\[PSG.8�ibe"1�2�f�L%��A����`)H��%T1H�S�1�!� �(�$r��J����#��B`����n��I���y�Ӟ������'��u/X�k�jbgQHA�/{�;�����?k��·kt��GQte��b�o�j��u���m���h��p�J�.ݰF7�n�=�+Dt-,z�����Գ�Q��ϋ��<B�M�'��0��t�9Y�[�' �F���r�ɿ=��V�����~¥B�r��"u��6����%�p���x�4[�0Mۄ����F�7����B�_��G�dx!���īZG&l�A>(�5�DB��� 0t?�\�ݬ�e�_c�' "�� ��f�B�;]L���ڜ!gr���9�]{j�R_8qHHHD&L�!��FV0lf��G��ܸ+P�)E������nvE/�w�v�f+?Y�9�Qs�$O�|8�i�Qx�m,�U�����ϗ%�;�������@����N'�Sͪ��&㈮z��7�	�?�S/��1��_L�4�|�L�:%���'�ʇ�m����������$�l�\��D���.)|Mܠ��C���َw �{�y���h@��'�ۯ,KV�W�ZW�������xR��~�1���� ��2`Z%@�kX��Sخ	�V�P	���:�޾�}w��9�ьA���Bp��	Ϧ ���Qg	�KsZ��T�\�V$�-����nQ�~,&wF�rJӻ�p�䋐ƐK��Xn�k>=k���7�UGWvT��{�3��BT�*'��}�؅�Sw�߽$>_�o7����������8b%ؽ��>�][]�z���2� Tu(
\ݖb�tZ�ݾx}Y���x�T��K��V'Gmu�@ݥ�{�Auʹ�_�<�3�9�!��p�a�t�V�)v~��W�������[u�C���[�T���j���!��NA��կ�>�w��Ĳe2{���Fظ���c���PP�����k�+�܃m����C_�7�a��v�Zss�;U[��N��S�)����`���HR#0S��;Qv��U��of��C�f�jS��q[o�3W�Z�O�A{��y0lPA�q���j�����9��ּ����Tl�`�GMx3)�"�	�L���DՆ�3�7��^�n	<�CUF��Ff����G��-�w�`A�Y� ���*�D�y6d�N?й6O�T�g���\�o?�QbS����.V@����Z�o>�����<z�ǣ��fs�Q�e��lAϗyr�F"-p�qUTA�T�;z6��!+��^E�٥"�U�x�	mIq� i��Is����.~��Ħ��`)��u���'d�d�H�|�git�Fbh���"��t�?���b`�	�A!��5�~Ĩx��|���f�L�Υ@%���P�aq�D�0�=eB���2���8������QSc����d��b'W=d�Z��x"#�y5���PK   � ~X��_8
  3
  /   images/57489f55-55cc-4ea4-8258-f1cf3d9c722d.png3
���PNG

   IHDR   d   .   �!�^   	pHYs  �  ��iTS   tEXtSoftware www.inkscape.org��<  	�IDATx��\klW>3���?�vR�ql7M���aBih 	�F4��hS���H�

�U���u� ��[�(!IqS�R�j�4&�;i�:[�w׻���|wv���cg/�u�I��uw����{�w�4`H�b濙%�k
�ٟn�N�W�éR6���KCCC�v�����$I��$���|�aM�<p�@ʿ�Al@2vPq�	�L��᠎�jii���2ڲe�,��,��=�}��7�~�o�.>��~��Cs���\AY�)�1::J�XL�c+���b����0E�Q\n`6�?a�Z̜	[w�\��4�
�"���(JB��|>��}\��y���y�j�̝�h��t1 ��������X��rrr�6�������i��̏2�j����ee��UUUTQQ!���A�Xyyy
�(>ȧIp�bA� Q�������w�gQdvk޴��;�oN�G9��9c�ڲ��1��Ջ�x��^E�2�� vݫ���vH*�Y3J#
��Sv�y�F���|
!HT��By,�|�{�1J��i�D��O1ױuT�y|բ��j^ՈcwH�V���RJ��@.i'Iי ��L*H��ͤ�wyh��3�PN�������v�j�**b$}�O���#� 0ہ�����TZZJK�.�lc� �������137~��	�Ht٫ju��+�Q%���3�|��a[Hz�$������Vjnna�֭[iѢE��OD�@�c������������Gn�;�>�Z*�B�QP���u��r¯�����cتjz�p���OИ]�/3_3��_�����0��3�K7!ǝ�xvb4O`η�3��"��V|ְ�y1Q9n�O4M�.]ҷ
�"�"��0�M7� 1�a�$������h�8.o6j�0m�{�<y7P���'�lo&c��Y3���#�1����9,b �:Dzd���drG6� ��O7j��41NG"#�L��Z�4>:zs���H�̤�1�!e�?�>�|��b\�)��{|k����8v�#
`�:��ac.$a1�1Ě����2_$}�`��[�P
b��LwWf!�a	��T.m&� c�
��b��(�1TU�'��nJ#YɎ@" ����I�������@�������7m!�8�m�9XFB�|�]�{�r|����5 �h���T��)�!_���b!L��_YYI۶m�ˮ�>����0�}�k���N�ec>�l�J��'_M�ҫV]UN��������~����w���"d����.^�H�+J� 4���Lit��g�-[�M�����A!�����g�v�|����vwM�I�i��)~�9��(+$g]�k&��+W��,)�U!Z� �"����療��D6`%��� 񋵩��O~�܉?z��G���X ��$)\��˺�|�k �������^��h�����C�O0	h3�w�*w�o�N��p�7�Ap��W>L���p��OJ͗Y_t�|����Q޾ig��o�7=!����?�)z ���ڵ�x �or�Oix��a���YN'k�厰�dG؋��\�ѣGi͚5�v�Zۑ�b	�+ H�����-̳�=��)�03qc�AQT�V�Y# Az{{EZ�������S���&-A���I�:YǬa��|��i��	igS�l�1�Ng��|�t�YA,�Ę���Ux�՜G�W����kMY{� v��g?G��g��lG�$��q��MI&K����l�anX�g\%�*c>�\�<��,�F�)D9����R/��]���q�6� �q���"�W��3_���K��9tn��w�F����6�m�K�u-����`��XS�JЩ���1B�G��������n%w���HԈ����{TRT�R��DR�����yqu�0�G�%^�1k�9���+�]��z��8�̿zK,�~�oJ�EXz_گ���JJ�"�d��@�ŋu�m��wۘv�iqa }|q>�t�q?q��v?�_^�����>0Ԑb���Ⳑ�]�z5����e%Is QN2�3�ļ/Fr�S�_�i YEx�~���2��,c�,� �t�b�!�!������"�z��5Q"&Ǥ��b������ҵ@΀�,��&����s�GI�X�e�(��܈��+A��X�`d���&�dd�/�L{�rB��bx����DVbĳ�R��Ф��7���Q�$eOrр񢧵1,���/��%%%�����l�̉ �P��������K�:���6���Z@�c��.
��=Â��g���O/Y��������]�Q�E�\��46�]̇������6k0'Q�}
�Y�v�+W>��Y�h�U��7���\��� ^��z�ϝ:uj!��9s&�����d�?�`]�ḣ��k��(�ǌ�Qbd����-�Ik�S�l�C��%�KX���Й��%vO�g<���شc�aM�a�}�=�
�7    IEND�B`�PK   � ~X�IM��  � /   images/86917e2b-5e70-481a-b4c7-aed39e2d087b.pngt�P�M�ED�~�t>��J��"(�= �	�C("�T���B%� ]�=U:�C�Pn�����Ν;���{��s����Gm͗tԬ�  �N�� �
	 ��s�*��!k��u�Wƞ ������r�}  n�ʋgz~ikxH,;1}�p�'���tn)E�EG;��ſm�3��ͦ�+m���0�΢��d�T�O�B���Țq�8n5���t����!1w��?�#��M��έ=��ݟm����gv�CLŻ�32֋J�։4���VV֋� ! l��!m��)_��.�[��]α�S >]O`�_~(BiJl#r��lI�.� �`֗�0W�a��?ư���+OϽ{Q�����1\��yQ�鉄Lc��l~�}�(	=>\8�(��z画~'w?pt&eHCwQ��xJ���'��XHP�F	sI[�ܛTN��n�e_>̎�8iHLv;��+f3�W���i�tU����\� ��L�o�"pUMI��Ol���@Y���;#o�s��Ōحj8���.aS����G�Yײ���6���)�*f�r��`��������_Z��#�a\x�;���������n<��㛪�k��k@a�����v��@��Dy�]d��PUrֻ�����bJ�/���>����k��c=��BV�V���?�N�=g���#�:�|.ƍR���P�t����B$��9EҾv<�4$�On����â�gP�ֈ��U��o줼�ْ֙���W��� Yr�
��U��2�߂DUͿyv��L "�H��+��P�J��.>Bm&���N���&��ff��c�a\V\}w��<��A�����|}",0��K*2�����k滠4��M��7V�E�A�b���W��CH)amR&R����B	���M���3[<(Y�z1]Ǜ���F�,����\R[���J6���2�&T��,��n�]��%`n�w�4fB\�}4G��7۔�+.g�����k��;�˳��!�W���mQ`5���ϟv�f��kTB!�̄�	��Z�QS�e�~�s��8�����e,�3���"�=�G�;����C���1�\��3���7�i@@M�M�	>w��k�or�X�K�0a��-/iB�Kt�	�%ai�J��W� 俗��W��;kTY�<����H�T�g�[��VS<Zeֈ֓*]|q�F
�����������obE�|W�"�wD�Ԙǒ�+�=5{�n$��Y��{7hl���ͺ�-z�N?��3��?�ܰN+H��`i<y(�y��^�R���"�±_?�w9�M+���g�2���Åg x�����ٙ΋v��������k����l�eD]r0�i����z�2���}�&���]�k��zw8[�~�DRa�K022*���M.��:����S|R|�]%��x��8۔UJ�&���(�W�����]���A������
�	���"ͧ_{���m��{�	b��\��999c�$K���vsf��@śN�nX��c	q����U� <�m��S���������FG��ة��iҌ#օ�q>������q���xT�0��SQ����Sc��YԔ����'��ƭ^�8>N��-�rF�_;�F�)?o@|�ڴ�h{S����w�(�.͠�T��񒕀ُ����_߈_�`��?#�#��z}�V/�/b��Z4�A�%�`��OĉU�Z#A]=���Qe(��A{�� {�nu@<����莮v"��2�Kr�x䱶������Ӝ8yoε��V9(L&W�k�M�r&�D�t�����TW�&�"M{w�\v� ������*��Qm<����2�g�i���wS�G N�[{:Ϻ>�yu%N��k���N��V����F]nI��^Ҹ���3ׯ��~R98�l2)���"�u������_%�����˞8�2@hkԒb%ĳ���_$_�yD�\���/(��K����]N��`��M��o_������X�#���k���G�.E�;�Vʠ 3+G���<;m/H�!{�P��I-+�Wפ%k*e�wih��-���	B��;خc�jD���}����?ybbշ��깠"K�u�J54����-��7hpѫ'�Z�ʘ1�ԑp˦�)�T�&+u�/�F�y��
������7����%H���ތ#sD���rC��\�\u&��'�|�����m�?����[����t��kN�f�9%&&z˝&�V�x4i��bT�^����^����>���:w����?��!/K��j8P���㿹?�&b��=u��	[�<=]��T�᳻(�.��n�YA�x9�{��a���,��Rā��/��|ҏ�˻�+�k;O/��|'U���</��h�J��o��Q�Z���B�f��b΍�A�NfF*�4�f����Ir"ݹF��F�.tX�R�>�1(M�J6�QE?^܏����<b>�]-��)���պ4�%9Y�ʤ��?�߾\�4��a[w%�UD��q�)+S�z�~k_9?�I<��a����G��Jᖻ&��q$���L݂�_ªx_f�BW��"��7���i���*��OX�K�,��M����f�3%�#-�:��3�������B�a��Z0�P%&e��8���Q���h�d(ۗ3��2���#�F��#�[:�El~���e�o���L�G����2���+Cp�zP,�>�^u��e����,�Ӽsݭ�X��.3?���Mx\�~������թy���5��]���F܈��U}-Is9;d���I���q��B n>���7:c)�P=�e��_�
�?v�B��K�<�w�����L�M{EN�� +FF%��=h��Ν�]�tN����<r�y���gha<�We������/�ؙ�^n�~&��t��m|,��pך0�[*�zeZ,Јj����ږ�0������`���G��Wx5x
�9�DO�}/�ǥ�S�2~��Sm�����F^��`dpc6���7�m���F��ݘ�j";�£�#��3�֩�oa{�.�|)fe?�I���7�m,�}��,z1�U�i�ľ�����!Kjo-'�j���)�{0�/W1Ex�ğ��}Z璱�^�F�|�����U�,`0�7:33#���E���f��x�T����nKU��т.��!X2ܻ����%�ť����?-� m<x���k��6dJ��!T(�.������u.##=�cXG��A"(W+�F[[ M�����;�����U��/��P�ØWI@"
��#�ݝ\5]���1���#�^65�XZr?u"�OOO	y�^3�W���yZ֚��6+���T��ZT.�Y��X����Xsã��o0�yD7�Ƶ�,��bXȠ�kx�tT̖�<�Qe����]�5��/�U��ܾIr`6JJV��P��s��Hu����k�$���[�
�s��$n�_��r��!^�$	�F"�#r]�V��Jl;���|�2j��zy���]ש��#1�b�!w�3�B��j����븫.%��d�S[��;�����u_��٩�t�'ߚ�4������;���2��^4߇��=Wk�A�Z��4��K�$�<;�&%W�eR��3���>+�@J���SL8 0�0Q�%������Z��L���V��o�9���>Cw[���OOT}E� �I|��p�u1���Z��}5�\�7��y��_0�3��l���Kf�TK�)�����3�����g��ݱ+�'OV�S�����.��QS4!,\����
\�������,��9gʡ�G�͋�?|~��ZT1?�x��=�`xnLKni�<>dbpz����B����{a�[����d�Cv��(��f�O�'�1�؛Ҿ���-ҿ��F�E�/��/��?hU;���QvBP���'=��|���X;���v��I49��J>��d��c<�ݖ0gRgv Cs9���m�E"�������R��Y��-�[�~�/AԒ;��A���~Z|��� 5�[��<HWT�����Dv!�Q]l�_2�?z�=�W�Mu>���4z2��b��元U����g�T�/�X��_��G�˚L���_�ƪf��=˖d]�o�\��?%\B6ʅ�E�@ �$vp0q�g'���?�N�L  ɸ�-��?,j�����P�o��k��QTj�\���'���\]XX��L5@�+�R���u8��/B긋����$G��͚�a�������ԟM=�:�G��Y6�{��.�~N�nd� h��?���҆3r�Ռ���y�LJ�b&}R'«S,����yH��duõD�ń`�l�����!���A��I��)���ߚ���q��@����	IdR����\�-o������y�]Ҟ�zE��Yb��*l���|G��*!=�A�8G��7}�y")`��<���Ɉ�,$�IB.@�
�z�>�:��u��a������w��ﻲMS`ك�l�\M��Kt>G�hŹӼ�"�x� ��ʵ�qbvd�rJ�����żu�hٺ-2�{����	&c�����_���c�cAT@��Q��|e��?y)���憽+������!������b���U���IaȚڑ�9+��E4-��Z\��z�]�E�(E�-i8�r�7�)�+|f���F��^�
\�Ԕ׏�yJ2{�C[���g��-6 ";���s27�;�Xs7xS��[�[�h��O��j���J>��R�'4���dzs��bAomqV�H���ǆm~�ǌX��ӓ)�ceBT+)uS{��ۤ�{	�}�ʱ[kr��f�i�x�cڂ"C(�`3��Iqx�y�%=
Zrh|�ED�����)��o�)���=}�Qr4�ҚSh�T��5�qu�^kF]�H�������6݃+�w͹&W[ME[-�q��s��`��X���܏3Ԋ �}Rn75�7�W#$�8�	;�z�%U�����JO��v��[A�g��]��	���4��l&|(-yɎΐ���'�ޟ�e��*�K�B}d���K(������������q��z6�X�Xv�!����b������İa@O�_`7,`|WϐT���t։�!
)�4V�d���£�>��ߜ��u؃u�	���
��*��X%_uz����KWT2�.�G���f�"��9��.1�COR��z"n���#�����ɕ&����f �Fۀ폠X~8������K��2Tp�y������c]h���n�ʬK5���5=�7����x����1E3�(
�b��]�3�B����B|�N�e�����VRώ{$��h6��!3�:��f���3d�C3�*V9�)���e�Хp���Q�g�>gux	��e'�Dc�An.�����o��~5���.G�a�����/�:�S3
\��	) 3l��]2j?j�H�ُ��XZ]�2xV}�:�=3�b@���	^!�W4�
�˞5#�5��u�����N�!��%^R�ׇ�¹P;@қ�����ۨ���1ͩ���ƾ���JSZJf*	VLI���a�Ѱ��q�J�)_��������C`�\���otú��ho(��#"��n�Jt��T^&��+7ƾ�n���$t����&ER/�>�HO�\�Eh0��淟UI(�I�=��c^[Ð��Dw�{[T!��bk�d�F'��Y`���_5�ҡ����H�"q&a��4�,[�0�a*0��2�htϓ8 �l��������z)¿���K�#辢6��ݚ���.ݜ�+����ևup?��*!�E�R�ˇ�W]��ee���M��{��5�,���3�s���3�[$��8��%�߱�g�5${\��'<��0'Bhel���1���W����L��Cږ�s�����~t�~"_28="W^�k�j×�o���ع$��s��%}�P��/+,�h4�Y�Y$&���� Fn����I]�n:���,-�x4]R�W�5����_�^R����fי}'o6	@D����R�m���y�<�dI?����Ax^Ĕ���i�D�N���|���Jޝ�~�?�/绉U�Vf3I�ݡ^���N!,�yWVo��͖u�N�/v#EA12O�Py-��Z�<�Wb�?ڷ�T�N~������kgD�a��{w�).�������9��E���f��7H��o�R�ݲzt�U��)�ƽ�J�"�������&h1�����O��l���i��Fo����
�{>���ť����X1Z�O��Y�цE����\yΓ�w̰��&.� ��G&�K��ث�@M���bB)]��E0����3f=좓x�,6!ˮu=_��dZgU�s��}���~D�`/ �O�u7J�&pV̊9
�zS�i1cnkf��WU�Y�wt��f=(!999���X먨(�)����i	�zj5�ͩ2�m�t�F�Q�Q�AS�;�斿�A���~���z/ַ�ʻ�1��)J�=vb������Qtp���gq���߾i]m��|��Le��)�TO��ݽ2V�'��~���퍛`��Ŏ�p
��6��3%�yZm��&��u5a^�3H�pZ�L1;*ڻ�Z�������gt�k����n����y˜3��W=���Q�d�^h�!x�����9XA8�$g��S
�adw��m�p�dw�Cy9t�dȥv�T|(i?�3zf�4��KtAW�_���F��B뽏p�G��X_��Ί�F���]������]-�&����\���ҋ��ME>U��Q�`bx.�#��._�$�Q?�ԨC�H�`��zi���za/�7?�ߨ���<2��)��>󊐡A�{��	./��Գ;"����s?A�܌��͌% �ïfntgʷ q��ϟyZz���N����L=��́A��R�e�!6x��ax	C�H������n���K��j
ds&��'�nb����NSa���[�B��䝶���B,�з߯���h���A�Q���d�Q���Z� �̊o�E�|��?��GD��e��Ų�scY���*e�i��ʑ�5�~=���)������Ň��^d��%L���S�^X�]�"�>������0�i*�R��X�h<mG�+5�����uՊA�B'���+̈��Z��$rt˒9Mf��i�ɕ$����]�i��4�H]&L �]R�c��w���d�&qI���2�@U0^�
�yA5�0aF�,��Cn-�w�#g�l
��Z��L�R8����;��T�>�"3�M޶2�����Y7���wwqI��Af���
���f�Enʹ�3`�J�͵�]G�8�HBs��a:��_��_����I*��uO�<��!a�-َ�A�FB����W�q���3:ۯΐ���v3����
�J<��� ��u4�c��	�Q?�,5d�PEHt<|�����*)��Mq���3��ҵa+%+��w��3�=�r�Q���N&!Y9��o�ƾ����5�e|��.��rf�]Yl̻�	k��o��gV�M�սg�Ş�&�(p�fXI��3��  �6!���[��,A�O���G���	��l-���Q��8�v�*iD��ҷ��]:�~��0h�$f���FqCPЬ���.�E�}��YH=D��7����+����|��'��UN��0��˘>B��g�!jyz�jk�{A���QkqĜ�����
�����T������88��ZpHE����1?�����@zU��-r쟛eu4&�\�jF$8�������b�ī��x�k.�Q�E9�y�-ε��<�	l�ϙ�Q�Y��KCƋ!A��7?��� �j�p��,,"޻Sgt�5u�w�LIT,P�P�u�T(��/��c:
�gqEj��֊�����Rr�9�D��|�r��FF{Fp��!MUE���
&)B���W�YG<��cx���q�wYX��2�;3��m\�QmY���b����+�y4dq��3�"�f�e^.�aAX`>
.���g�L�6p�Dh���m�q������^\o��� �s,�EW�=#��K�`(S�b$��2�Bv��VW��n,�����p��Q~����xg��ƴ�T��+��zۃ?Ͽ��(  j�/�r����h�&xC����\y��%��8X�f��+k�H�͇��-�ܘ8��?�R˝��xD�6Km��te>�|�m�T�Dr��?�|1��w3�4�;c���n،"ո���\���	�U��ĕ�>$r��^�&'�<��"֜2��N�G�|֐T������w3F����w����l2s/͇�M���}�'S�79�)�1oi4�i̔o�ۤ@�[�U6�Q�KI�$ܘC+���� w5!\^R�"m�$K�=��:`YY&�����Q�*[���J�8�͉O��T����>Χ,.�ppY6g�ӛͅ�R���B�	l����Br�8>�wR{���(��6���v<�x���H��"_��l � ���"�����֒�|��'p,b�P��D~b_�5��"�=m)��gh�ܪ�1���\^�(�X|f ��t�ʸu�ΊZ�d��a��=�9 }�M:�8��8,���:��8. A�Sg�u�Vuu�Z)�/��u�g�~BekLW��&$����.����kՙ�Ř�̦�H<@�E�S��9���b��l�����A�'�F$��Q�M@��M!X�rt��!}��x&֦���6����+V?�띣/�j{��Ѩ`SQ�g�B�<8(�n_C�d��oe�����Jy��b��3C���Օ�ޅ����mc���45�(p�S�r���κ��4��z��VB�>�����r�r��H�Ԃ.M��������Z$��p�3�H"���%nD�x}��sa�:T��ۻ,��<!��j���&�%��tvvu�z��Ĥa{/���G�-%hRi4�9�s������1�'	��k+J�,�ܩ���*�I�+�:��+i�� ���Ͽ�j�?���k�#�p��R��&s�>�.�l~�=#E��M�vk	��g�X���WL��|VzLE���`�ׄ�ce���#&����i�19od�dUԆG���Uڔ{�L ,��F����^����-��coY���+1�
|��6��A��'q����~��������Ay�֖�Q����҉7�=d��`���h}�wz����Je��>�M3��X_��!'\�c��x�N���E�Ɔ(����wJ�N��)��8�t��vH�Ը��U�}���[ٗ�T��h���	GM��(�	�1�X*Ze!����[[s�i�
�QV.9���?iʂ�� O*��[:|��=DE1���
�	���!��Ϣ>�ۣՂ�+�º��ӛ������v���B�n�u}�%�?`�Xֻq�����i�P	�c���ս<V�܎��ʠ��$x������Od=�S�K���q�Ay�3)89���u��U��?�yO_u	P���;���q�FxeF�N�Ȼ�lb���h����x��I�ܑӇ�KΝ�OW�cU����u6���T��5B/M�V\���e��}��M���i�	}�G;cL�%$0�1��V]X>\�A����o_KP/"�{�ퟎ�%�t�o�mG�9����(v�v/q=t�j[�ˠ�xJlQ��|��ٮ��k�d�9�~�����@��'�/�=�?'S���|gVfo{q���# �d(�H<=��~�V8��u��h�%���Tk��������'����ϑԫ��ň��v�:W�-�}��=~�A�;�aT�"��_��#P#~rdj
;4����FJ���Փ�t)�m�teZ3akl ���'�/�G��;H��}�Ѐ��H���(UF���K>���ŏ.Ԕsu����]1/ž��$[�����A�F�ݳ�����q6F̤����u<�Đ�3`�2_���P��h�3��
 lsõۢۯ���+�f3[1�����x��ČyL���?`�sx�,���$v�erg�l'�$ˈv����[��+D*�6�\�p�KA�c��򯜁�߶�=�S�1�P��w�( �r�K?1Ì�0�o�ū�D�ӟ��}}W�ژG����y������� u�jŻA8���jߙ�NJ���z]�'}����mj�c���颉����s�D&��͎����X/��.=��A]���׶ݳ��w���d�&�c��#�]ȶ�1��<M����o������1�-h&��ۻ�3$���f������2��7��η���pI�9��Zl�E\�����i��KAxp����%��Qw�qE���|*cfZY�k
n``�
^W���@��3�2����&#k����%�Ϩ(����B��KљK���"��B,.n���\娆����c���޹��m1��9ssJ|ͣGZ�������<��N��a���0�.��avz��^#�����ݘ��gdOt'?c��!�H��p��@!@���G��錄ڵb������ۉ��~�l�����Cc��b��
��ӯ쓛��	�v:BqYo�$_���لM���l��'91��u�=[�+���J����{F�(��愂�)�,�Z���/2�(�4�V�	]SX5�f�e����9��EJd�K�S����.���9�*�!�T�:ι}�DX���k�����=��屚!=F]Ї���v|����zv�K ��2D/��� (ة���-���8��yrM��A�r�J7Xʳ���LL*(���ڿ���v9��- �������;�)S?�����/��?�7���q��������"l�@1�� %]�3鷩Xxٙu;�x���>��)��%��l�[.��IQ�E'��������A\	ԗTR쎤 ���ۗ+����\��{����������YZ��5<Sڊ4s�=����^�'���Џ#98f���.|k"VЀ�ZCs��`7zy�"��d2����*��7���ͪR��C����V�I"\�kQ���˩�5L��"�����v^puw��c����&^7�]����.��"\8��o甪u� �������;[�\�cwoeO�{�?�$75aA���q�n4E8���7��u����^�_���Q�$&v�����^.�4�.w������	��B@���ڴf��+�Ϫ0]�9�@�P�
�l�̉�s�ʟ�����n������]���ȕK(�B����>�!�y�w��6!x�8B�{C�,�Z���j��/�W���W-',����"�:��ȼ]쁂*����G�=�{�*�2�?w��b\�3e��^z�#O�o�y���&q�+�%M����gq��W�"]�WW�2P�HF�)��(���1�f�U$X����6��e�Cc#��x��g�������D��*9�����ۼ��ɼlil(qRTrxi�H����<��_7��!�nV�rrT '�Z|#ь<���_�C���V4]���;��Q5�e?A\	��85+ҵ�l�dۊշVp�W���]���ف9����	aX��S�q�	�r���a@@ �#I�;X��ܗ�=Vͣw���r��*��ߑ� ����ܩ����o�ig�*��[�X�5���1�1�I!�Ͻ�*�nt���T��w�u�Kz��T!���G.dͩ�˛�&,T���E��{r.���5��`����1z�l��"wЧ����7g�Iߘ���GC$��̈́�ֵzK�sSG�s3۴�ӧ߯�M��Wn�� �oR2��N�{���&����i�1��L�o=���^i��=@�Z*⎮&P޴���lsK3w���^5uRW@�i�+�hs��|��$]�m���ɂ�>M�"�9�U�U��ֺF�;�p(�*y�!/"B��f���!^0`�m/|9:�W��8i��5�A/��P��l(�rOku)t?���4!�i�HϱiHC
Zc({�sb������F�+čGA�M��y.������}N"�$+��,����:�t����ְ��n��{p��$e@��0eq;���>�j*�F������P� ��A��
��(E�v�+��G���\�?��=n��2�<<4�B��O�N�o%��t�#O)�ޢ^F(������Dd8�=j��s��3����m�c^�6Ͽ�`3��&5]��㫆O��]lqU���M����g��c1@�_�/°�8�5�*�d����M ��0�O\@z�����O$�2�T�V�SΓYKHc䲬����3����=x��6ZN�9�=�ʘ������(�E�R�'�fOE̵�d����\-6Լ���%����6��휀�6�l�ؓ��α�s�GV��7������J}�㯐����Ϛ�=c���S�{:��$���`�|�Y�>v�=� ���ª���ιo�#��n��斫�SBLa��"u�����?N�<��!&C��O��z��dTI�B+��w��W2�jŁ!g-�^}ԫ�
F؛Q
��=���6�K.�0+�*g�;���'�<�f�>�K �7&��!:i�3�K$8G�����(s�I���+��)9h���򯆦��_ ~��&���p'��r��*�g8vn�KR�y6x�j�;�������U�M����.1�nƇ��y�����V뷮�0{x��9撒��rWc2�?m�1B���ۗ��ub�a,� 8���\X �I{\�k#zKU
`���Q�fX�?���o}�^�B���O�@i�sA���MA<���#�W:��=��f���"�mu|r�T䝄���c�{ބn\�*�zE4?����\n�r�5��^m�z������`7�4Dި{g�"���������4����vKy7�FC�N�>s�<ב�*[�H�ɣ�G޻xhXw8�5�naY��ԾŔl��g�fR��{�B*����p]8��vc0�c�I�s�8��%�fG�[⪤6��fi�TJ(?<o�1۷{S���c;S��Z�o��x��2wQd��t��ӏ̯nG�u���E8R3풤�=��ܸ���١�P�n���ц�`i��ԸyfϢà��CxO����ؕT�*�P�D�
NC	|f6ɷ�QR"�
M�`Wg����<����fv���h'}WmMW�Պ����*+�gɐS��B�F��z�}0���v�t����z�o���l��M9��^�����%���������E?����e�g�����6��Z|}�X����3zNQY��vS�a�S������sMGUģ����-������֭������VS똣Mi��A���z	YY6�oPh���Ij@݋���K�����{���{=� 곆	�������fr��;|>�����sm��Q���V����,.	k�ג�%�̩h@��PS?�R���/䀬p_�ؼ%�[�}CԱ�W�N]�)W�"���©��YB�!{��Z �^,:��*㻮W��G��E���LA��<�B��B�ϠUF�WN�NX�z��BUy��]���ƨ\(bբ��T�[�Н�	[��9���[e�cͳ���9=-�FȖ��,C��Iţ�:���qI�g�< ni�L�~�Y�w�y��ʘ�~}��K�R�柁����|�F�y�OU`�aA�fH�A[���	���b���Ծ=���(����m���K��K�g�q~fM���)\�r$
.a������$��ӹyɲ���+M�m=��P.R_U�[�a���v3�է�Fm���T����"x��7����W��&o*���G�zx�o�S�h뽜^8,Ƃ-b�8Y�0�a��H�\;e��lF対��iV�>&��Ÿ��;1���@�?i�+�9���>��#���7h�%-2�[8����SgSk��W���U�Ee��nd�5=B�X䲂Œ�!t�HR�Vab�EI	={X)�-�#<��V�xFC�ڤ=a�E?�X2H��;u��wY���tv����8��!g�˙��Us!���R�OG2U��m�T����u��j�VLƑNX����)/ܧ"��aI���%���^�_ʜRG�1�ʵ�t����=K�"U��h�B�oZ5�6:d���J &-��KF��H�X��ZLY/I%��稱"WA�Ī �G�FQ�I�@z�|�ƔX�üK����>
H!��#��˒�A5�0w� de�?X�:�2v�úueE5��`�R��O���_jFF�Ǐe8��Ԗ�u�b���A���#��z�4ޡZ7"uq��]�l2��#�G�9�W�6d��E�-=�K�TV>��/Ԋn�ܞ��"�#"S���t�����y1��g�k�f�&:��:�H�����h�B��R��w���cg��f|���7?2YQS�\��no7(6z� ��3..R��u�z9g�o�:��Z�<1�|���̱WaGo4�e�P��KN`ro�wC`ɨ��tW�#�J�
T�jC(��
�lH�:݃�uN���L��5GQ/��v���6��{mN�	��EG���;	�ŕ�P���֬TM��U����2Yp	�phiu���Vݩ�GS��Q	�td0"����_����I�xP?d����[��t'�6+E͔�U -��l��2	�ˡ��[�'�'S��了!�}w�/�w�t�����m_��"_����7� 3Y��� !���ʑ�r#P=�~�B�'p��P��/[�	�l��FNM���|)��Y�Uױ�灐�jtr��<@7t+S�Jl2��T�.�z#^}���wsL��O�Z'�8���s�`���<�x�շ羡�UD��V"_~�ʺ:~ӡ��6�I��.�T�'U���\b��b��X�5E��E��ӓ֖xw�jz۵l�0�Á����������,T��TT� m���+@�����E׌2��d��ISW��1>��KKރ*�^��6����h��+V�R�$�p�Q�1d�9�)��)� A)��냁VS���ဇ}��'}��K��^t�g�"t?�w��
�5���#�;��/����Y�@V����{��L�@�NR���u���������W������\�_����y�^��xt��"v�
 �]���/��}��ywl�>*���us��"��f^hi�2�n��5����~%���m��+����;��'.��2 ��^�b�`U�jC{���<��<�<�-�3�ⶵ;I[��u;���C�����Y��e))A2���Li��-<C��ky��b0�9�/Ä)k��vꞱ���'�C� ��YA	�o=��A+h��lK�@"ָaO�j�r�PBg+V�-���? [�w�N�g�� 2c��z�L"��8ӣz<֙B��P����g����#Z=ߩ�]]]�� ��H���K5�&��S�n�g���g���YQ�9ʣն��F��1��tnʰ���.��R��!�\u{��D�KK��-��IЀ5�B�L�������&ʣ2�T���)L2���x�@G��L�?Ϸ�﹐�qXI'tt*-�t��]����wq��*��n��2��d�+��1�%���� �������Â�󼵷@Z`��B���ު����H8�����7t���/eR����T���|�>*��!�W��$�x�@��M��&�4Ҕ痒�[�������g���A'���Ru���2@f�g����^�#dSðS�%W�am�<�
n������ m��b?��|�]�_���{��=���e�����I�V[;��W�8�D��&�e�[-���T�Css���y��G��>6���G�I�B]�]�������/�n��~��Y�¢�h�E�7y� �'Js>���}{U>xٓ-B[*�>�6Z
���D��L��`9�K8�8��&%�Kv���{H�2�l B=3>@.
�M��?ww���. }�I0Y���Ń������Xv~y��l��Ez�j� �9��1-_��ش���K�_��p洯nd�2�#&ί��k��S����ps/�`P��ϩ�E
�\u��3��4�<W����I��gڌ��JU���*!6U�r�K���;t�[T� �]�A%3d(���:���7�w�6{�	Ts�82ݟ�^��7"?�G������X�]p�U�P�<�
؃������2|䘶���k���A�������#Y���ӓ��'�h��ʶGX�g�hHi���d�T��q�(R�W��@W���w�}��?X@��s����bǎ4����vk�է(4	�3����>��/!��O)C�w?���^)�pv9�QT��X�Vg:����H�agqW�UC���)��$�=������R��IE�L��E'���8B��	�D��LjF����1���?-o��>�a�]���"-c� Q��&a7a�,9�H������E=���I� ���͹G�Qc=?���ߙ��O���E�=�Jb�29����h�-,3��<�6�N@!0�Wa�OJuo�5l�d%]��n4��C������|��w�B�8�@�29�mDN\;�������3'�H�*S	�		���d!�2��rk;'�F���!`�/-����^,ϟE@���
�"��[�7+���[%@:/��)L��0s�O�ݧ�,)�b��z�r� ����vi��A�f��Ɨ��ᶉ�\�p����� +Gӵ���9���J� g����X�i%T/��.ɘ���(�?�����f��n��������ao����OJ��B��.��%;yG%�1ٳ�c�k(%$�:$ی}��6D��}7�R��Xg��o�?���|�����������u���:�\#i*WlW�W�ΐ=�Kp��K��:�A+�k�2O�`��Ce�9�_wl�]L
̥^��on��q�f)��J���ԑ)@Od��c��}z�S�F=͑�X���r��s�@m /Ņ�2����ъa�1�F�(�$�V_*�SH������U�987T��A�7�ʋ �5ٽ��K�(*�3%!.��w�d�������ꆝv�����MO�Q�`��Bb�i�M#M����ktfۏke�b�	􄸷�3����=-���i��^u)������_���ǟ�����_��p�ݲ,1ЀM6B���嶱v���gG���^�,��<����`L�3�Y��%��ÎO^>|�K��'�s(�P�������HA,��qZ�-�|m��"�K�b}�\ �M�����	�V�����Ϗ@�A��~���Fn�y<����t���Dk��&bz�$	���!�X��Yi-FZ��R�a���J�
ms���noyt�At��L������,��V�߃������֖_��zv��-9t�g>�<�cr�x�t?R���J�,Ò7l��a �a�c��
�aN�3�0��
��_�j"�V��s�j���D�av�F�J�#;�����n�Rn��k��{���\�� ]��Tζ��W-�w����.}�(�u���6x�,��`�U���w��_�>�$���ΛtD�S����~�t�Y�G�uKԍC��<�uW��d�,]��\��Ϲl�b�������s^$���@�7+�:uMM��f^ߛi�7��1s�_�_�;�Uu�����gb��� /#qyS#ϴj���:����ZS������0���L��L^����Ҩi�YC�n��l�Z���\�nz��އ������,G�^�n�ؒW�0�lC���Ք�c�^��v0��$Ǖ�{6�^��o��F+���xǵ_���A���� ��_΄ e�=O1]�w[��y�QC�O�l�&�_0,)��`Zm�97cW	���o�4�����c�V��L;��_�7��͸{T���f1��?h��<��S���)�WeI!ۢ3+D�R�61�ѷ+����7�/�,����)���'�;�� ����̕P��z�����_s��mY)ȭj={7��Wߣ�N{�����a��'�4��OU�ú�6�L��QQ��3��`�z���`��"�-r����k:�8
F��c�.L�O^*X��u�f�8O�b�[fǓ�r�^Lb2|�ogLx��VIڀ%;��<�rN3�"P���m��O� �x�ZQ��);<OѦ��H�<���S��]�>W���fQ�r�`^�=��N���|Ԁx�ς%V\���cM����'�K�ݢ��f��,����S��t��B�>p�ǻm���~�S]-;&W���DgeЧd&yt^?��������"�g7	�W1��{���z�F$ai��H3����
c351���\�f�������H��þM������kM]�G��Mj�v�Kb�G��8�Zo̻�a���".�U2���yw�MF�Y��^�o�;3�����偛e���bJQAyY���&/M��?�s�؟-�k�S�j�}�r$M�����r�W�p����Q9��}�HM����=�z� LD��*�-��`o?����2����<-MV�{�������z���A�u���I6=yw�z���)�� F3O�(�&||�/)P&�����j���F���,��+�L��}���}�hP�yO� ���d�d�qDo��  ɾ�m�&7ӑI�%.�S�������8m�vN뗨%�./�VT;!��b:�ӻ-fM;c��ȑʜ�ͼ�Ѡ�]�b���pyA��,�����g������ii��L����Δ�p$�?�t8A!���fyw�Lz�����y��Ȼ��H�P��� ��s�J��¿�)�@��ğQ2�MݘZ¶ފ,s`�=g�5��"�� c�*�:��*I���"\A�--,T	����c�L�f>���*9;������Ҹ�y��,N�̷2�� B����)�,N���~S���4�����ʳc�v޶��,t��� N�������U����mjz����ޮ9��[����$�����c���އ�;�4��9���&b��gHf����o���N/�p�Ҿ��i͹�.n�������ԫ<�v������F����&nT�bl�����'G�kQ�϶XW NT
������ެ�'b���\L
�TƄ��X�~�<X�qr���v�����Q�Ą���F<��& *��/S�AMJ���0&٤�k,�T%����cW	�8�&����QU��m�<�85@!�������.�.���D�&<A���~4��I:��˶z�oA�)��>wo�	�r����({SeI͓�>v|U�*�ýa�O��]37w`;���i�������?o� �+@;�îo\��#���*{�}�����f���L�^Gz���-��I7�Q���=p�
#{r�~U��4Ihr��\���^�~�u��Ʌ��w���u~~_�Q�s(���}��M^R��-6?j�\8��8Kƭ@���>:�UeG{:6譙��(.����2Oo�9Ø� �_�`��s�z+g噑�����e��&yQ�c��M����� ��XO%�z��t�ɭ1�E����}S1U��Akd"�������U~7�?��R� _s���n*z�Dא]����si��Z�eZ�y�@�����������e*�/zȉu@;�<��Jh����>u;�ཷ���Ӕ�A��x��rי O��E8�S�z�5��ϱ�K��[��5����p���X�b�}غ���{��5V0�ݎ��sF����u~_��r�eN�h���F��vW�#�d�Ŏ�_>��B��� -���޳.��k�0.&�(q�5��oQα�/����A1�����.Tğ[O��Ĭj|�F?֝����^�?�_��ۖ�<�-���ƫ�%�;k�P%�0�V��9e��"��T�L�8ƴ�4�S�yz�8���!��9oȷS��Ci$�6��{F{��n?�Dy6�A�I�5���"�3��!9m�s$.g����"���-O�1S_��1  �ɼ�+8��|��ѿ��@5�nX̛�NS���p�A�j�7�n��&U��K[�IN��z����[7S��Ÿ��f
wxj���&�W���ɵ����=���~W��B��L`qW�1�u^��̸g*���;���L���N��e����!�~�������e�\%㎼���nv�|�+�_��܁�2KVje~rܮ�-��k���c�O���i0ip�?-~��i  <��97�S�n�����1�tJMƴ0A����؛��6��%�0H��C}�#��f�0M�r�?�n�ؙ�sě}���J�c�����+��b;1� �{?����� g�VF(�<�Xި�&���%�-?�.J�	3 ĸ��vh���z슌X�W�y[�ϪR���U� g�]|����fA��	�.�z6�e[�l=Sa��<���e���3����W�'��$�ׯľRs�D]j�>k#2Zk�T����}�� ���\��3~w��[F��Go��)V��[d1�oo2d��ĈptXr��I�� �$���.�^��{���`z��ڸ*�ePբ_��l�~�x	r�7���h�������� f@&f��i��(>�ĸ�&`�b��ը��lT�cN���yx3��h�A*ǹ�_����I�ݖ����	1�{��01f����t�V%�p���n���\痋���h��[�F<�ty��M7�x-@J/ܼ�{hbUr���o<,����Z2��H2%t
�CeK�7Qw��]��~��&�q­���>C�L��R�|�Y?��{���b�돋���٘�5��>V^/�͑��i�G��M��]���ظ�:�����WoԺ�m@��	�e\^����Kz�܉oɞ��{{K����c�P�9���\���ȉ5�����lb0��GE:j`��?i5+�^��9��wd0)K
��~�&'q>�o��y��F� �_n~�!���M���ה�f���>p&Q狗��P��Mj|T|�?߯n�'�?I;�n��s�f,�ٕິ�Dj�~;?;7�C��*8u>�E��D�����=�B�:O� ��u	Y��H����OuO<NI����҄c�e@;��Ϭdߢ�D�'vrk|nڬo�v��O��^��$!l06FR5�����"#Mȁ�� c?b���	�;�#E��x�=(aa㑤Pqqi�����ȼ,M[^���$҄zU�Q7�Հو38��1�=�4�x��	q:W��ieD�a���εU�/�{����W��N+ߖj-?�ҁ�ؿ6�"�;V����U?��dWvt�
L�1�I�)B�����8r�_�ȬA����mzg]]]/9��O���_���]��Pa��V�ƨ_v�O��ɗE�2�7m��7R�0#�؊���F3 �?*�g�����Z���-��ˬ��l����9�����!9�ӛ�g.����Ο���;a^���G)�'D�@)L"��?��0�=�.1c��G�vԕʾ�� ��Ƈۖ�b|~��6=R5�}��K�;��43:�M�ۏd�����s7Y. @t�Q�y��u��goe+
;5M�X�$әZ�0���B��V�z��-����;fR�<\��3�Y�`ͭHT�����Sr\5�t��+�<�KԸ4�>��I2-��z�9\l�H�tz����Ѿ#�Z�j��[A���1��j}[Jc�LT���į9��w<�/B"6���[������Q��m�6u���X�d
��������4�ٟ�L	��)�l�6S���y�ޑ����zɑi�NR���罏�+�Z~D�.zE�R7j��n��I�~s��g�EcU��a��K Q\{31*�1��&�Ɂe|�{�	��Z���j���^��@4 ��d���1T��0kwD�1�\G�h�v�*�,����O`�t_��9�T�d�8�X�]w e+Nai��p;���wE6iw��O��h�:F��p*lU���"�}?��X^]�s�~`�M��߆c|����:�UMV�`n�.>�y�~3��dB=�'����<���� g�-Q��'J��u��{�ؐ?�Cg=����v';׍�B�j�H���(�i�E��[#8?E���O�Z��9�Fc�t��y�Pa6�1T�_z�׏�/=:t�8�|?Q�57L��P��y�pR�3LN���T�E��B��ş�]FO-g�6#~Tܨ��tF\�t;GuC��h��"$=�5��6��SSO%�"-��t���N/K��Q*Pk�V,E��=xaÖ9"��t�vΒ]�G�n�c�c��]��X+O���P�i��34r�j�}[�M�Vp��2-Zz
�w�*�h`V<݃6rT>�y%���7鈁i�g��r��lM8��������)�r���8j���-��7��V����j��m�V`�G0���W��@���*��=|��ތ�x���j&a�IM��PnW��wQ�CꖊC-�\~���'���~*��1Z�j���&L��1�vS�� �v�~q��)/����nm� ]ǌ��p��4bW���n�m�#�?��d�'WURkdm���TS�
?E3�h�] �D%h���ܽu������
Ʉ'�OϽ5�$-��ob��~�`���Ǉ�aL�J������=��?ˋs��������uwyr(��J��C�l�)h:�k<�Q���P>FbK�^���ƩI���A���-R�Z�n�x-�s̎
���]�	"j��t�2�� q��N/ �|�����#y��mi~���>�	\��UvG6?�˛����9 ��1��v[������C�,�5�L��W��'A����+���hn��}�G/ʮ~�>��'���q�1_�YR��Fk��   V��mD�1�!Ş)�Ũs+\�z�YY(����Oп�a�{'`�Q ��m�7s�#�����T��:�̣]w�$I��>�کv̈I���p��T||Z��h{S���@���R�$�3W26p<�>��[
�x����q�a�t���.æA�T������^Ml�����|b��&����jTOKe�r1��o�
�^�vŎ_��߆&�,��"�n����)�`�~�y�<��"������ڒ���!���ꬹ�4���#��W����Q=���+Mn��$�O0�o�]}e�]2.'� ?ggg�n}C�8��W���X�Y�!����W5�L",����!�� |�٣�KN�T��ѩ��6����؉��N��+��G ��v**G32��f��׮����8Ώ����i���&~�^��;��vE�7��ZI�t�3a۴��HP�!f�σc�ʐ{�У��F�M���������t�u��[1H9�!�O�& �4�`��}���?����I)��Bp7�Yʢ���#�ת��؉V�t�Y���G��w�e�%׈��u��[���
}��k*~�0jķ���Zw��V �b,;�7s@���磿2�-��)@�����⚪֤ޏy�M��$ªg~b����\|8�K^vC�� 3�w
)I% -SԹ\D�Ŕx�O� ���P��Rn(�������h�sg	w��\�V�F:�QT�HB;��NNHo�}�Z&�M��[ �d�p�����N1����%��o���VBe�g��R�C��<\�y���D�(�Y��}|�+ֆ�Yݷ>_.�m�'k��vՌ*�+�.��t�{�nZ�G���?3x'}�U[���L�E��5H�Drr�2�����@���X�zy��6�<��ל4S94�I��9�=����#`sPض����@��K��)�ئQ'��	�§�N��6>��[���`}ѱ����^�V�����6����Q@���o��7��y�rk�
y�r�9`���,�=� �c�{}�3BJmp��;MPvIy"�I���Z%�7���"�L�[��6�]=<ț��R\s3�@m�����$��Ag�}�]��>��Hd�}�6���� ٟ�<}&����.�xYJ�_{k�!��Ӌ��31�׹k�g	���o����E�D 5��[0G�Θ��l�S�h;�\�VeƈL�K�����N��yP���{�,=0�gK����, QE��(��[=�����]��0���7x%�,FTT\=�@>>��\.H�)�Cp}=%' �����h�ľ����"[]��G���Z�}�,M[!J0�&"�5�4-g
�/���z
�˞B��� �I��ɕ"$NŁ�ʃ����\fnz^�v�嫙�oΫv���}�٩(�s�P2^�ٿ2����{��ջ���o��|8{٩#z�ŋ��������I�^���X�d$�+�h�F^+g/4��^pF���j|�����X!
U�?��-	��LZ<yM(��*��e`������Ķ�)`�:+�'-�V���mMLL��=<<neU�4���]$�d:9}^{Sl�DPZy3� o��/�+�~�	p�:��4�Y�]Su��r�ys���I8Y�i�fQ��\�`)r��C-X�=U��;�7|O���M��$ ���>hfO��2��E� ��U�/-3sT���_����V:fw9���ٝ(���x"�"�1�'��n� R����~��I�[~=(������cff���1P^ڻi�8��7FY�^g�(�m�F��dĈ��D���K�߁�qTd:�s�&x����u"ؼ'�U�����ws�x�t�'����A��0RtG���Ɛ%�������J�6�[t��t��>�
��D�~���H���i�g��gg�u��F�������A.�ZT��ӿ���(��
�e�>)k���V�n4L�W�{�hk]a���NA�겆���uh����%F_�0��:,���4ޛ��o�,�r.6	Lqz�y�ީ� �!Y��sUOe�s25=������P��-M�+�\N�����������n��}��?p����iC�d1�����d�t�	����B@�|��m#uuu���?N�窿ƻ�qƋ@��z����&0|E=� �l�������X����ͷ7X3~�U�M~W�\����yn�4׆��LI�!Z=��e�9
*<��E�P�z{�yF�ز�(���/A� 21�	���&���N�c�0���K��eML(����������y�*�%�����dT����1�B(�� �5}�p�-�e�A�`[�c寅����at��C�kjk=�&���UU��L����b8�g���@r�K�o�{��몯�>D�YH�'<(�q�=����^~M������U��E�/�g�<�h���ݙ�ܴ[
�BS�\V���\��s�IO��}�����^��ع����k<�o&JѴ�����U���U������~�qO5��-�`¡�B�(Y�g"�e���x�X�\�iz��Tp�>+@1�`�3���Y��Ƴ��j�h�Q�s[G �oJB��z���n�����yA>u���?ƌ���t/�l|���9`��z�JPI�w�x�󍪢>�K��)����Ѿs5�/L^:�~g���ݞC,t���5o�(�.�h���$$��� �����Ì�"��yT0�ٽjF)ȰK;��D��T�!* 7�q��R@��KG9/^,KII9Iv�r�6�<c��#�f-y�Y�W]% qб1C�\c�:}zls�����gf�;t|��z���^^^�,�tȌ�����h��@}ȃ��>�wۉq�����7��)����=�Y_��h����F��׶����yz���ـ���ɀ��B�dOUT�[yRH���v�Q�Ea���N{9؟���#6��e����6|�2 �S�z��T3j+t���塟m��Pq6S;:@�ΣU�GS�Ffn�
��-<2�LR��'��T��w��詩��Q�Z۫J�	��(�����������*M$n��cjϽ�G_�gh����Q�5;����bO�C�y�#�t�臡�+���^Jy�(����$��������_\{�v�$�����U/hb7�}�|x���2�������'1?���f����uDJͰϗ���fUˤ7�&峣=+��N�R��!c�{���xē1ğ�5���i��ѧ�nC��z�mgŇy�����5�v��tI����Ww$��_����)���t��?��^�0�T�9��kc�ӄ�l��|���g̦�� l�قA�>�����x�}`�s���������AJj��ȳ�v��n)daxz`��4MwW�r����$�n�[&@r��a��7��
���� ���9��&d��B)�M��ɾ�8�ώ	C�ZS)cc\7ve�ןg��q��7�.vv������򷗖��k��e�!E�Ω߹�s�j����g��kHEhP�aX�k�-��&w��?
>:�	�<�m컷�wJ�Q�ݨ��ny��kך�LM����nn�@&$p5?�͛U��(��@
<B����vy���\�nπh��ji��lE Qi0�0Dy�4��V��D��ρ�ٞO��0� V�pQ�~��h�����X��? �����/eo1�w��!�6^+��k
ս+6��N�d)�aMr��M
�X�޹�h�2=C�i;��Z��p z��vI2H�{��uO�\��!S�|���0�옃߯��w��H���8*�h�|�6~�X\���GE��aT}�Cu-Pͅ��JV�a��f�6���kb|F��Hʬ�>�iG,	ڤX�'=��Y5�&8�Pzm[2l�;ܶ�NF���2�a\s��~z�y�B�|.TV־���P�X���P��XAS7��>�n �vNx~�a��ݠ��y�X'<�02�A���A�p0������ey�)Q�|E�W^���ATޡ���has��n�r�TŐD�X�1Ec���k�j6�Vq����SCL�\=Yt���h�y��y5C'��X��g
���-m?2]�������Ct�6�SGyB�	q����O޷H�a����%� �W�A� �/\(��bA�Vh�eʃ���I�z��ax1i.��k�kۍ�nh��'J9�O�]0�?�q�ٴ�+)sy����*��ƹ��w�j"��ȉ�����1Nx	��/�)�
���jVr;jɋ���%KȂk(cB֠]������G w�q�����$�m�ݜ�����Ъ��Y�S_�!��Ň�G�{��P�NŜffA+��@�L�`��8zr���,�3�����O�����w2	�I[d��3E��)�D� |A��|�٨T�א��kp�>P)�3
U3���dg�m12�d�o�z�dG��k���ő��㟉W�C=>�IX �����M`�ǆE�R�
������,T��f,�ؙ
&׬�cFH���̶&��G5

�j���/� ������z��ޝ�ü�)��vv�P���Ȏn��`�����ߐ��+t黱B���eI�e�D���<��=[5z..9�L�A,��G�[���$x�:;�a���M�`R�:b-[��Lt��W�u4b��L�:�\vz���o�=9A����N���F������="az2hr��k|'��)�?����+�N��*����<r�pM'���;�`�$ҩ̤��a�^T�����bD��|�og���#�����ȡ���N>3|��3Qƽ��'?�l^�*�8�4�� ����9�\�c�8��*ٖ7x���d�����#Jv�M�ȿ�6PD�@%��v�?R~�C���^"d��|����]"���iK�ML<��E����c��A5�����G��vݟ�/2��B���^6��� �,������r��x\1b�M���cVυ�ռ�WM�P<��Q+�m�n=��v�t�� ���~�����|ƍ�����eL���cq7�#UH���~U�m,�㫍��!���M��Y�0	�r�X��7��,�ch��~�;�Hy��A���M��a�B�xWb���ұ�/Q��u^�޳&�I��h��`zG�o�m�7Kx����N3�F�W�����
�$~.)�~�+k�9����c-
��o����ڳ��� �`���2��l��Ğ��=��w]ZYҕ� �$R�{ Tō��;d�����i�]QN���^�L �1���
guqt� ��vm>,}�>�5C���w���9<�]3ܹ��6	��^��z#����kb}4����5\"�\>)���_��04�Y��]ܜZ����
��������-�T�h{���&�c���� 	��)��r.��,Ɍ_`X���p�6}��g1!�p8+�h~q~�Pn��G�e�R$������o�]�؀�U���G�\�z(��� ����L�S��%�s.3����~|�?:Ϭ����/6F�����57�	^q<~���yk�ZM%L��UǉB�v�@y����~c*&��a%�r)l���n�*�UbS&r���;bXc��c''�ba��P�}�W|�߂��a�̀�]���Z�kw�i=�,Pf����?�����=s�\��/���NK�@,yPa��^�I�3��5���r;C�Uכ����bX�Se���R�mv�j�ߛ�[��řSk������Ģ�R{�z��b�dO�]E����5�v>��:M�}.�qP{����0��Ă��Ǥ�% J����� <"
��}U?Y�\�b58��q���Q�C(U��3o�~wW�����慑=���~
��n��_-U�O�H�7sC�E��~șM�qD���	
eF2.��y�p�Jr��/�)���/�+�>�d�A�?QI�
%w��Xy)�:�o$���A��8�s�����6���v�ޞ�u9�:[:�n��̸��c��%
҇��3�M�F�~��8�����	�/R������k��H�bVxr�[[?�@7ϰ�zn,%��{��j�ڈ��j�"/�Tv�o�%����e~BSAu�n<|0V,&�RPd�d�K�=q�����l�l�ئ�|��
�LLh�>~N͞�2��cv�o`̶֙�JCo]��~������Gp����
� �+~�q�Ο�^��V��n�x<~��I��b�<�#;���5�6))�h㞼�aV�C̾X����f����C�ׯ_M!�/�K����y��pԐ�S0�?�Q	���/A@��J�	BN���{:�<5����*����+�K򍿹x�pag����o[5�
r|���rS��>/�q�������@�H���c�q<Z����'���ǯ���yo���R]E��>�<�\�p�6?z[���T��!%Ssk����5m������	�5I�zhn���Urr���9����J)u��a�z���iG��D>i��,����s�ߺI��`�x��/K�))��;��ID����D����m��|�4Y��={?��?r=洸�(�Z�!�V�аp���Z���i���nw�`�p�����O��(d�g�"jd5�;�_�84�08�a{ol�
%e�8��Uw�Ƥ�Y��;���7�6�m���O���͍LG-l%;Kuk}T�+��
��Ɨ:�.��N9����]�ƀJ���������D��-�:S�=��FF��K�w��`(b�^��Z�;��;2��fB�#��:D�i��p��nU]Zz��S 
���bbb�MU� �S�\ۛ��B�J��lXnk��^ y��,9&j���9 ���@U4H���u�|�p�<Wʣ���AW��=h+_-�bov�P���c!���7��������z�ˎ�L�ۘ5�^	j	�/�����k��c�f.��N�O8R��kΥt�I�֨ۑ�g�A��M?Ɲ.i�I�?�ň�A�a�.���t^�����%��t�az���B-h	�C����_U�Tu*)cv�v�Zḋ'�~wNu�ݖ���*�dk�-�7g��Ԡ� ��h�ۀ[⇗�R�r�5�(y�c�lk�������K�]vo$����n(�S�&qRSe꩝��:�ȡm�<G�2Lk�w�_���WUTTƟd�*�FM/���6���'7 ��G�\`7*���Qg��҂b��V�a�4�p� �=۱�J��QW��-�-�s�9����T=�Z�ݵ읝���M��*-��p����A��Uz[���Aנ��4$n���:�,呋Yٍ�Թf�oO��QČN��Ի��(|#8g�ylUVh����ƚV�T�!}t����n��]��Op�����gee��%������!����~��>���n-����%��0�������	�<�X1�z|	9��}���Cq	����lq�k�M��9���#ʮ�įCH"���.�>u�����`��EV���SH���p����m���2���&�ƫ��L�e�c)��]��+Q��2k�}����������.I�L������^�~FXXG7�,����k͈��p��h��i����l;��s���\���B^�&~�?�"����?|�"���+W�"b�¨���s
�j72d� .���g�F�/x�W�+�#d�٣����Q���ю�9���iJ��\8�o��	}�fjH�>��A6���J}p#p�>�y<z�5Z �if����a��DI���x��ʘ\�f�t��3ߥ������B���3�O�3����W|(���^ipG�t�T�|y,eK��=�PE�^h�]/$�&F2��@����s$�Ӄ-�\�/�W�-*�=$g,�f��
-Ɗ��P����D��T�sDZ�ax�C�L'�7����ʞ^y'�}`�돑�.�}�j��i?��
�8'����D��a��'k�|��tGVvy�E ם�ƶY �`L����I(�ь�P���Q �v�_�&�-�j&��רapb[���~��D~���}V��N�@w�0�z�8��Uhm�o@QW�l�Hm��q���?�F��#��'Qp��Z<(�p���z��^	We�w�.B�~��9�V�8�T�w_v�Xﻹ􌈕5�.���6g���~�P
��sK��F�-�>��ρ��~��t��֏/H��� o�Cw䴦�T{f}�@.3�m������h��Ғ^E��DV�o-cbJ�k<ږg@�x���`ƍ�}i���˪խ�6jЁ}�(��\a/,��p��鷛�����z�\g�z�y�o�Ӈ��~ !B��g���r$�qyˠ��M�@���xf I�����39���͍�/����	�R�@�� ������s�Bb%
�T��An�OV��u��J �Mx�|j,����AE�aU�,wuv��M0����5��6��A�]�8�h����Q�W��ey�f`�m1��GA(�o�=���N�(ڪ����i�< ����s�z�ss��1��x	���������5� �_���vc	�'cd"�E䋿�1���>$9k�H��U�����R|�*5hi��Z,���p���ަq"(�f����p)���i�����X3���a}�j�D��R�ӆ�Ө�\��Ɨn2�!6�2Z�/2�rh+����<֍�bs�
��5�}8���ӍB���9�����ڱ&�B;D��}
K~2{����i�y������hZW��1cT:t ���2�*�s]���g������O���'PJ��"*�k�v++������0�P#MMM}2�����x�L$�{�s�����5$J�q�%&LZ�08��yb��8-qw(����16��/�W��(���a_2y�'�RҌ����0���Ws6�r���5���ncz�O#+�KH1g�+z��H(���W"�7{ngJ���?(y�- 6�t0u7@��F^��{���P���o�Alw3Z�T�~��n���C�*	�4��4 ���[��u���j��=E�m�9e�T�aT>k��z��7�}�(9T(���&^v���z	��׭�~oz5!9�����*CG����>rV��1>0/�ի�E���D�P8"g����_��1�:}���ݻYOD9nף�!%В�-|�(h&�ٯ}�E�3퉭����������˷�����չa �{a�B�+L ���V����H<�o1@N�&6;%J��U�̃�����t�?�/���'ZKJ����7��M�8��s)���
3�Eu��f���Ń�2�	����8��@��)I"\����ڝ�s՘+k�ZC��Uƣx-���{7��D�-�H6F� ��]9�n/���ވP��ZbFI�����$�~�I�=Jx%8��S�>-�CLn�D�nd�^���Q;�L�X�v�W�5�3��w�oy���)��H4 �i�~�6�a>�
:Iz�AXv�.�qw`W�G/�)QW-X} Q6���oEC�����n�iff���J�~���|k��\8y���Y��L2�z���wD��V��D��/�> 2���y��tXW�q[g��i��E�bJ������P,��[Rmʴ��A�a#�i�CQQ��rI/x���p����ST��}1 𧨧��Cܗ��.����{���ԏ�}}��>��a�?!P���{;4����p�F]L���w%w-h���{��`?"##p��ǟ�$�6�d�d-�$�ppH�\���yH����X�~-L�|�94��DsOO�:T޲	$@Rԋ��믨K��=�#� �L��S7I�_E�5����#)�������1���%6����
iy�B��Aȹ!)+{i�QSi�{-� �[)g���x~5y����H2�M�=�%F�F�.�ǜH����P3+�_���EH�$�-�鲩�B���f�P��HG�xwk?>74v(�RgA�q��C�@s��\��%_�ӿ��\o8b����������#��HEi�c.��;W��R�;wg�w���<��(���-.a����+Z�X'�ď�w������Q�e`>o��VG���@�d�o�7�2��к�?)ciFQM~J��yQ�� _�=ӌ�H�4�%��N�u����V�J(�3洷yth��p�;�s�-��FY��{��}��)�W�E:���\�]���jx*[�� N�����u��ԟ�@�n&��}ȝ޹������&yH��z�Z�����)�M���e}��|���q�e	1�X�+��Mb��^�<�8_%
��K�����
�uL�7l�p$�� <RrG�䫆�nUS�Mm���6�!c�c�mk�o% ;�y���O��-	�o�:e)�������7�����(�Lh�/����'}�0�h#�̇��*.%�-_b��-1,>���[L|ì��>e����Iס�E�F�[�3z�+㮹څ�v���p5RR7M yN�c+��H逅X\%��c/	��h7�a��wU]�#��F0��^LެA�����t�|�/�տ����ᄌ2�šf��Sм[K�h��r�dA����^1@�J�F �4tˈ8�ძ)�n����v�"��tr�4\�6i����B��K���œj`��g����v�!�ߴu�E��j8���l���C��K�=�PU�����c@	��3���+C^+!�<�}��ٜ�D���%�7�ON�hLكg�T*�;�MOMI�%!+���?.��Q��J ���R�Bw�(Y�Ĺ?�-�r�<��k�#��o��f�ع0cȾ �S�K��³�y����6�̑P��5���z���KX�	�zH����;�+&��,�_\z��.�R~�l���,�_yH�|�����4Ld�	�X�J� �jM�����X2�dx���`7=r�<p{k��;b�&�H�G�G.�/�\���k����ƛ�$IӴ<s��Tyc-=��/\��~��g�ʌl��K�Ӧ����(�5oB�^cL5�r���ǀ����+����Yz&�����#��|��a��@��?fuYE[���J��ؑ�ګ�L�5K[{ob��EK�BlboB"�����|�����"ו����\�q��.�Z-�W���LQ�[�,��>~r^̣����Xw�Dj�g�\�6B�����
9`֚D���K���ۡh?{���gx���r��,͋[��|q�z���"��s�2L�?�}�n],>��)�>�&鱐��7�z�a��r����"�uRꗠ6�����
�4G!p�5{�CD�m���,��ӵ�:��(>�X������GZ?	�iP�C-Q���犆^5�O�i�'�ɽ�PmS`�?�&�h�ٷ�ӱ�cx���F5!9-Ox�[#�ޓ�2�k��i��9 ���\���f�^i�F��0=.�~�l? ab�k$ �'3`��S텼�2����.�c���g��W8�}N�.�"1&I��h0LU%?�VK�^Ɯv�h��<�Y�2��]ﰣ&(��E	6��i�4<�G6���z|���0�b��B�f�6n3��`��|��KU8ը�	c���H�gF�^��1.���5|�%a�����E�N��=K}�a��VD}���Z�)D^ P51X]n�P4i������AȄx@�=�eqi��k4®f�"�P�C)��ΏE��$�%
L�U�}�z�Af����{��:��amQ"�=�VS�Ov��{\ױH2
��R�0�K$hM�	L���.P���{��p���C�ɘ��f%޻�c�{cC����C7�)7���C��<������;_�X���b&Kۏ���MSҠ��F&
�捥B����rk�|mt��^��>��x�?O�0x~�=��!�_j8�*X�f(#mA�����c��=.q��Yv+_f�e�����=��Z˾�u6_�&���3 ��M]'��N@�K��.E�[	�&�$Eu�2�2���R�J-7l�7��a��r̅3��\���N�y��w�y��o5�hn�S\�<�$����Ѽ�s�/�I�]T4�����|HM�ݤ��R._�2\\-�<䛐_�/䗃�{#��v��E}�j��ߐ�|��.�C��f9Jq}&LF��C�; #@���<۟������uO�}Yc�µ��rH��w�����To�o�@�(�`�#�lΕx��a����d{w�M?k�4�>Z벪�����0��rXn�?��Ee<*�k�u&臅䓫�T����7�Z������k���O�����Qɱ�n#*9[)V���3A$�]g�/���Yc�����G�3QA�G�#@F#���=�N8%_��1�k�/٪6���#��IH�y��'B�X&`h��K���m�m6!����5�O��|�w� it$��|��o�����A���:ﳗ��.�s`]��̷���hE�\;b��P=��1(z˞���-FO6�?�"�{c��������D*���.]646fL�-�x�M�ˇ;v��~��uz�ZA���8
��6��cE�kD�p
vV�q��H�$�!�'z�R�?6jRω)�,��1K�z�1�z��}�7��lֆ8�A��N&|*�m(w��X"ͣ�/Tlؕ5)��u����I�ƨ`ǵ!lȤk�Ž`�c�vU���o'�q���j�8V[��4�|�5)�zۣR E�ċe�~]�7�8NcB�iw_^��l��p�֧��Y�żv�pB�vuN('4�����90�H��]8l�;�
A#�o�{��A��4�js~��nq���K�"������Q�J2��}�!.GTF~7 �L�P槻Y��go?",q�`k3L�g7b��� �D�q_�x�V%:�oD�6��:�B3 kI����Q �K��B_Rڦl�;V�O�ةB����=�h_.�3�=$������n���Y/�ދ�,sW��E�3�6(��RP�ʟ��Q;�@��$���K|���X(C�����7v�|����C o�m��S���[�zWl�����CUEn�l�i�F�_�'wk��;�)~jjE���]��}UpU��vN�>�w�����H����(Xn5f^�[ԩC�-�z���h�:ܡnU��8/��{b�vs��T�ҭ�9(HJ����$xGѡ`�@1��<��-�&O�B�F��������q�����y�(+�vK��+D��J��U<Y��DBN?�&v��55���/F���!c���� ��Ec�M�iDS����<Qrh�Z��a������GO]W�~]�S��m|���,�^P�o�U�G�g�Ʌ���<?�������5��n� f)�7Q��1C<Q�f�0��t��-�^�6�ނ'k6GSfk��gz-o�5[D��U̲b|Ф4r)�3���{�R	�/��ܸ��w��r�B`��;=�p(�6�	�ޣcTLY�ku�2Z�_�<��=��h�׵~���ha��de�5d�B\\1��GI`vεeQ�󏩨o��x��!poI��1@��]b��^3��8a��4x��Z�����L-�ue����EU�������6i*rtndq���q�`w{?���̇l#�>��bAQ�7r|�vԟ�����8t�����i *���up�W�^�w/~�hp;�s�����E��D�<�Wl�w�����;\>��i�.qE�Ĝz�K���)����O&�Ӥ�:�|-2���e[�ޠ9�2�1�g�����"a�ޠ�2u%�Ύ�!�r���sj��0��^^��@<�R���|Z�y
��������\��s��R:�|��Ռj�Cd��l��d\,%j�u�x
_�$=�s[�Y�g�2W%���M�"���]zl��Ps35«*s/Y-��j'bTYF;�����:��7����j��@��K�:��A#y�;��B[B�W�;7'�5L>`��Am[�q�7�'�w���f�7��gAF��jw0�0S���E����P���4Za5|�g��2��Xw��o��� V�����-w.M����8?���g�b���}b��O1�Ǐ�N��K���K���}��~�s5ϫ)��UI�Q]���u ��1����n��[�6�.ܚ\~�j�Z�8�*r�<��g� B�>��A�.7�!>KÏN�$
��G������}��H-DV�G�J�4=�S�nY{�>���ﳧ����'M�a􆰷�^C�d_��%�W ��\�b�O���Xl�d�ޘ{���. ���d�c�Q#)^a�ibd�������7ɽi?Ԧ�C�@����9�@�h�x�O�s��J\��K_�ƍa�C���/zi���z����c�ө����WVW+>|���ie����mG����-
)ge�vH��H�2&&d��5�S���*#�ER���1T�e���h���+�Q�� #	甝WE�=���G&<����_u�I�{�t0Oo����!#�6ZcD����վ�����Q�^1��E}�W�1����:U�e
h�c�º�Ӎ��ueu���wZ᭦�S����$���3O��Y-��T9S?�[îak� ێV��Dv��e6Wʭ��;����k�˒B�3��6����$.wݽ#Qu��S4���$75��r�{����U�:_+&E��(����f~̸ۀ�ww���Z�΢�VW�����n��;����yyN�ڷ������`5%Y��W&���%�fj{�eA�O�ʇؚXtZ�-�Y4�d�WkV��8x���Z�Jm�mS����y���@U�٠�Kw�O���/qEJ�a4Z@�hs�l��h �<�yJ����K"��Bw�)��I�֖�f�ۊ��z���Q��$&��-��L�r�S{j���ZR��X9q��n"&�qGKP�������#���r<�H���,�j$��ׅ(j��.�U�8k�E MN$H���߅`n��ma�-ʼ熔F�3k.��wx���\de�)ڝ�ȎXf���/�L��$sz��S�pV�k�¬�qc���N�:b�l�����<���ݘ?�(h�u��s�`��������{FWI� ����+c��zHL���XG��F��<C�R�ȵ3h[Iϋ�_,l<e�4�_�9������-Q:���a||��K$5	��ۂ8u�z�B��xX����鷽�Mt�6���]�=�P�ﳞ��V���`���\��5�}QD��P�����IĞ��f�/���jM���q�i�k�F�����F����G�~�	F`wR�Uy��`�ȔLNZ���'�(�mi���7���y��G�p�����܋Q5¹�!����7�����*�pܿG���8�|8�(#pS*�[�l&��*^"�_� uBh>�R��o�\�w�7�j��+ĝ�Z� �t�g6z&��$�n�q�S�/B�������/�����!=��H��n'+~[g��"LY=���x�D�7��d#܈3l ]j1��R�4jM@0�k��ʍ���d+c(��ﭼ?="����O�:E?T�:���[9�Uv3�;AbE5�����_=R��C��]ЁUש��?K��^T* �WI*�S������__M���5<Yf�N�ŗ	잗4E3՚j���?�{��G�N�q�Τ%��Ɲ��:[	��wo]E�~tQ�������U�/������7�`#1'譜��t����X�՝��8$\d�G[�RK��y��~A��Ҩ�	�M,�4~ �ڰ1��tm,+8d���M�>#.��J��}<���b8���϶��cZ���d�J��jj�c��{�}�1U��A�*�ΝrI������`�n�����i�]Q���p�7���(�Rr���<� O��z<kj���og�?s��`�]_q�V�qqIH̎�5�����J�Nw�h�y�����t
���e�Ct�K���m�����cq)Ѭ��:Y��4���:>��@Vs�#�$�� ��@��obn�ܰ�7<Z�-�b	�au.y��9�`~��NȨ7��I��(��4�k+���r�wP?�����Mz�>����9T�yW����͌��3|�ڨ�b���������C�f�j���s�O�An��(na�P31���6?�M>8�ǵ��������hC��N�`&��t�d�`����|���&A�C*���5�7�k1�<�g<���65�������7�k��[�M����K���ui�ƻ�o��:'xh ҉����H\��絺���2�Q�*�8�U3E��A'�v��ߡ�6��6B�-I���)��9��8�X��q8�������t�;k����l|��7�ohn|y��������R�
�5!OTnm�<E7�c��:�E	�㯜µ��5^�b�U"��7 T�Z(F&�x�Ȋi��ebI>8
�/y���vA��*�	�O��¶�K��0��,�
Ė��M738�6  �`�=�b�[�����9/N� a��Rg^lA?Xt3/sʪ�c��ݿ�e"q5FF?����6:�'3'����:��z-�vf��t�q3��g\ e�w$5�k�8ڮ'��q뱇����Z+��i&l�8���O�$f���|���zl++ѽh~p8��� ���>YΔ����VW���9l�O��4/��
�}NLӤ�Ηn��#s��|d��ƍT��3/�� ���G�X%{�C&��lc�~��y����C]�py|�۴G�6�.ɒ�V+{n���NA�E�
� �`���|�^~8{Z�R��������0��3��R
�A�6���pW-E�'��\�b�~0Ԇ�8�n���Z>Z}4^��p5t����$�q��
�M����U0��J-�aJU�i�9�U��`����p�
�I�������}�v#p[�=z,��iק8����oB�����z߀?�B���ʟ&l���A<.�!�0��w*2t�(=��fj08��y�n4�EAe������$�O��捼�򝨉vb�4���*f�8��!J^��p#��)��'����" x���pe�Ğ��6��O���7�<(��rRTB{��;�a�Ǎw��$�~�X��oa��O냠��O�y���&���ĺ+���ib�E����,y뒧P�����f�e�j;�K5�Z鬴�d���deօg���{�^�Y�T�%�ѻ&����x�*���u�}��n��oSG�
�^'��=&Zs;�Oc8Ӹ�C��F� ��G(�{��f8�7��kxs@h1��wk�i@�5��d{��d�.;���GPص�W��6�� ��4�����R���G�[����ݕk�q�YT-ѥT��F�Y�$���5��ëF��r�i^�s9nsm�T?J�5�1��g�2I3�O�9⪾-A�H\��?��?�	�ؑ&BVO ������L����%�6QSRU����t��zR�:�K}�l�����=0�lnhӠ⋖�:�=/�ȶ�������ˆ[�t��Z/��d��/B?�o�	�̐�@�`�q��*U�BȄ�a���>au�3��d|�-��,�h��(P2�P��(�E��$�KUР��X˪lS��B���װ�H�]['дZ�Y���\0^+�bF��(H�A�7�&Z�Gc�}�t�yɐ�6مi�I�����+�������-?�N�괈�
�Jt�c|-��/p�z��Q.0k�B� ��~i�o8z�6��K�f�#���ۑ�R3-?��5��'/�u��y�V�Ք�<riYu'�ܼ�z%n�o�]�%��Q��%h��~��M��,ۻ�l�v�,z�
�Ū�_x�f�7P*�t��\�#��HA �k�K�����&���		ǳ���f�+I�n�ߟ ��%���dm-���v�����ï*1V�i���`�f��������h��@�޺0 �ٴ�W"�B��,��F���Ij�m���*UH�,6���>n���cAe�魼��B������9_֤T��lI�8� �H����ST�=�n�}��X`*xgQG���̷7i j��O�#]�}-�h�B�HEn��+�?7&����0�3���$�"�;d�O:H�&�|���3J��5K<����qԟ�:� g�/�2Wc�S�sX��NC�=��"�vG!�'��d�"�Gk�}�����XÔN�qe�}NiQ�Q�!+�ѳfH`'_^g$7vh@L0:,cd��^o��_:&���d}�&�S��� =��M�K&�ڠ|�Î��iq�,Ү'G�6�ؼ���7��E�X���H�m��fS���z$}}x�����jZK>z�F\\<Z���:yL������Ja ��i<1<8ɣ��h���-�u5Ё�Dn�	�6�IIr��^!�\!�˟�}���&�5��h��W��\�x��ˤ��A��=i��-��������oed�%�@gZ���*��_���+h����k�+]�y�=��`�ˡ�v�-���P/(֫=�)���o��.�'h��o��<��,a���-�o������#�_��\�ypO�	d
��/N�3P�0Ɣ�]������l>cx�q��2�����r���a��>9�R� �RHh���f�` .<�p����Ǹz��Q(�I�h����QAM��,�\>zN�b�@�v�-wY8 pܒ/XR,;��lx��3,��
~�>���ĥ�f�k��\9\��^���7�n�12ɇܸ����?�vY*��yMy�M=:9�\tc ?�1�d�����>�푝X�fsZiJ�
����ԝ�U���:;�a�嫡�.�09�)�m%�(�tx��?�d���C�CQ�RX\���x[�������\;�f��$��{�Z{�SP�ݸʆ ��|x�\�'�3m7vsT�FTxhJ�-n�%~�a/�\9�_i���if�[�_N��˟�� �W˛���@�}Χ���;����=�pcֆqy�C�1�}�$�aZ��<GC���7Y�ymF:��,x&�$��fj k���%��;�����n�1�b,�`�3*�QE�F^� S��z�H$"�����2>����g���b-����l�"p,z���>֦���:��;:u�Y��r�:��Gvz��#��П�]^Eo��Y��A�O���h��1%�����O�2�)Y�F"���,/@ bm�`����؄�;()�GM<�k۾�Y^6���h�eE6��qV������Ҍ/x��q�@�WGf$���U�h���~�s�4�	`w�����G�`�����p6�&��b�c1`V�h���ϱ[ҙO�^&�9��V�	��ܹ�:p�߬�IÅI��3�hDa�k��BQ"��Z�-o�`W���ԨW���:�?&mTr@Q�okF���w��
l4@fC�g�l�����6��e�i_��0O͸#�d��R�>A12f�q��Ք��R�D�8����䩣�D�J����V���
�CclT@]q!���F{�lđ	��n���֌ri �<�9t�V�B��j_P�nX�� ��ѵY��r��$l\�:�7�=��������+I0��+wl���ۦ��{��j��ҭ�!�0��)r�KvY� _�
�ѽp�ts`� <�]i�v׵������ҫdd�Yn�k��Am��S�2�/���ٯ��߅FysW4��}G�~��3��HŜ�pZ�����vu�/QP�
��@�����:Fi�h>��� ���=�5P�`>u����Y���ft��<zR#�O�2�8tL��y(J��y`����|hO t�6ٜ�V�ٱ�=a��"K@)Q�x���v>S)�^��3Sek"�8��5���R����\�B��{Ò��Pd����7�'���yyۓ�z�[;�Y|~�]�|��8���1��!�
�Ҩ3��MV��lw�^�3��sh[�y����`�'�l�5���؆��#X��-��2;恱��n��RyS�G��ּ�iȸ��u�l��R8���53��v^�Ϟ]y�(��(F����S����]39�Q��t��:Ąmm��� '�<�[�������<���U��v��H�ʼ�����Ν(���|ԭG3��zq55�q$޺Τ�Vg�w���2%�[�@[��Y�h%��uL���^�5k��Z�M��E�懽5K���C����$�b�g��ؾ��M������۱��zM��m���=�/��i|�v��DaJ:%�w�ꨉ�ZM˗�k0���}nޘ�"9���q��h7�1�U;#���|�&.�̘��k��.F�pV/��y�lȽQ���K�Wx�Y��x�櫉o���TY��x�{8M$�ϑ/[%G�u ����n6�d�5�����H�˟�9G�bv)v��]��:֒j��u�2��(�g�{����σ�Y���&�x�1���a��Т4��J�]Mh]>�zgW���hi~�CTh;3L��, '��p�qղ"��*90�SW�jd�Rb��;�#�/322x외]��Q�����Q�ҷq������Խ��ĉ�[<�=��L��U�T�R)�V
L��2~�)���B�و�\�44�(le�@6n��o;�Ub��ew�$��"b�Qjl1�C� �^2CS���L�p��	������X��&� ���r��?Ҽ{�c�`D�]�q�>=�r`����>9�)$������!��*�1BH]1|Ȕi�t��E[�>�.�	"�����-R�9'�	�)���0�]>� uI�9E��՘G;�:��LsFO��2J��Z>\мs� 4��,#""&d�0x������7����@vR!��@�7� g�y��bͩ�Y`�&�yxmNYU\�x.ǩ�U�������~;��Vԭ��T����>;ł�\Cc�8�PF�u�x�M���*AW�9��B|S}���z�+Z���.���r�f�wu��]�~��f�)�b��T�b=��F^d���=�{���U�`ү���	A�1D|@�*p���E��S�{�ָ���o�5������'�^�5Q���n��wXf޹�xa����Ӝ(P㻒+��xp�d@#�V�x��{;�-'oȓ�O~�sY�тء=�s�ۻ����+X:�HqZ��e�:��}_���F��k�dB��8�B�����6�9�#�A���Et�8A��0r��ʨǦ�dOHe��l��� ~j���s��K4j��G=	�\���;����SmkϏ,������n��\v�,b�����I'��J�>;��>�����՝�D¬m��۝��#�ή����qq� ��3Oy�����v;][d͹�ڢ?����wü��r���' h�վ���88�q���H/�f{��z�Q�0��ލ�*g�����/�b	�����r�\���}��^�ԧ�Z�W����ϊ~ҥ?���v��q���誔��G�.KL�@�b��>��n�x����gHct��L��a��1q�kV��J�j��޾~Z���_&fx9� �X;�\7X��z�V{�����tGN�$hY�>Ց^�����(}x��cM��N���rn�ݬ�,��=/zV4 (�<y��?����k�e��b�[�k�3�c�AW){�<�dZ�z=�n^��9�ɺ�%��4oo�l������k����3
4������'��*�C��\�?Ӗ�j��r�_����zw��3;�Al��r�=<$-��Po1�ėӒ5�g�w�� e����:��E)��&���
H����u�D�#�`��W�U�НS9SK�k�����P�C!��"w2�ފK�Zv���R
��z��_fv̾F�o(#i���]�1��xh�m��`����A^18]��W��`ژk�{���7�4��(��t��̴{��璟������%��gUA�_E�����?��8/i�sP����~��!5�"�L>�������REZd"�&����PEin��ߤ|�0Wld �>Fɪ�:��p�U1�kͧ��<�潏P}���&��~�$qе�~�U�� ��/t�_����޳�#n��k�5�N����F�\��\�#l�l�_���F����(/s��$��>|��$n��ݝ6���+.�_[�L��&��`5>shT�
(T�}b�\>����q"[� ��2�_$!&ƈu��WS��H��_NF���/�+QmlC�]3��U��h���7�R��w��ws���
T�SW�tJ��!6���Z�9G����1&��r��ŋ�i$���+��3A���ެ;1���]�Cm�<�3*�(pX���b�yq^D�:/�����-U��l�Z����ej�Kc��n�|��F˧ȇ��ؓ�B_�lNk�3�Dūb��u����C�@�1W���;��o�3�Ѯ�4�V7"_SDY���!�J��Cm�����b������S�V�������q'��g�nU�I�2A�d _�a���뎽�.��M���%Q�g��p����?#&������¿�����]���X�^a����b'I�$'s'�oSP��(���B�"2��*:�|ݶ*Ǟw��ܼ�Y�3���Ԇ?�0ӌu���i�	)k�I�}r���z�h��Z�ZsZ��F�s�r_x���v�%���S����1w| w�޹>�Z�r��}� Co$�j6@��;h)�����r�`�Z��$$h: BسO�.�R��R�!(�=GK��Vq�'����q�\�b�꛼���7�T����_���V44z�Ѩ���V����(�{V�O�mcQ�LѶ����	]����~�'�8���_{>_��J[��6���Mjy���GGs��o�&+��?���-}I����;�
ʟaǰ9�ձ�����KT'�#�=d�ڏ�TD��ƤVx!�?���&��9Tu����;B��ɸA��䢟$^���O����dr���/P�q��UI�2Ϲڛ���h�%F�}4��MU�X"8b`v� >j����d����|�B����xM�2:��n�Ql �>eӎ|P4�����Ǧ�/wY_*g�c�]4)����؛w%Ը4@�߻�iߍ'P"	�o��R�/�2�Dc�r{_q�1^��g�M=�^+���P,{�ra�V���	g��b��`�C�K6NA�0P�nk���J�~�$���u_jL��o�Öp���zk�;N��}��.�e�������ܸ`hd@ؙ�üjs��ro|53����xGHl�0�*���5Q�<���+4���F������ep^��x4�ݽ�MM�Ɍ����+��p)���8��if��*d�[_Y�P\1��d��D=��$W�Z�[G���[�Ř���U
ͫW�j�V.����2���C2v{�z;6��s7�-&P2�贿xS6�TbV<oӲ8}5���&���Χ[&ϛ7K����,�y��J���o�R�z\_OF�����sbw�P)�ٔ��N������+�_��/w���5c����5�)�� ��F鞙�ʝ������2}lD��ÐS����P߷[��Äw�?d(~Ƹ��y~X���ce���PKi�`}��
E�>��"D���Q��.��n�)�2e�;�E���)Lj�����2�� �	)���q|�·�W}>�������y�'g,�[q2���v�@�n�`�!?���+ȎOU�w[�����U�#�vqyLP놓����8f�f+���I�ur��J ��5�`���
0&fb��r�`#wE{2�Cy���cń��?�j]HzN˭����������J�.���@��z�z���a���l �XQS	�y�25]o�l}��î�8�L�@����0�'��mT�g���(gv�o�!I�-7��b��CI|���\�s������h���{GOϑ��ǕIPߊ��4�'���8��d�l���:�X ��i׌ǋn��K��h�!��Ρ�r��'��r8��J)�#ȶ���(�6֤����s��Ub��nQ�������ޚ_Š��NJ���8H���/c�ХP�ye�[�Ӏ��J���}�Шֹ�;��˸ⅉǺZ���rOl��� E8IuY���e�zΏ�B���bi��[���y_��]u���}�{��m�=�d,��;�vz��C��o��;O*a*_����f��7��[vdؽ#k3�{�M�S�\:H�Fw�E2(��j�Q�B>��ɓr�^�?z�ܩ=&�]�Iٔ��~������5�r�Dh�F�zĪ�F2��{�!6��F�����	�^��_*��}k��9��Nu��T\O�prl؋�s��~�0������ُT�%��KorS�֜֠���
��D�ӬvUU챷�kC�I�A7��T����k	�,�$��@�4��Ж1=0�P^��3��@����e����(d����-f�śdd�w�Cb�����ߑ�K��v�O�I�I��c��Å<c�\�=�(0�'o��0�8�m>�)Rcv�����K\�������su
����n�@��!�::�f�IT��c�Q�g)K�z�xO��*"<��p�ݹޛ�����l���\�ZF_8�������T
L�[MR�ZJr��;����H�̦�e��"��a�݊�ؐ�!j�2��a/�_ ���K��N������'$�֚'�ڪ��IՕW���L5���/��v�sƁ��~�{T?��|Ϳ�X�Ʊ��#���s���;BמF�w�9V�D�U��N�̕���=�Ew+���B��˨ڥܤ�.��U�4�(4nkk�b�6�+���N��`V�
�$=Q��j�?�!�q3t��������&U W��y��.�+P)�/�F�ҋ����+>��X1�	/����jT�KF�	���#�{���ħ�z�������Wٓ�]�T�������oI~���ȥ2i\�h=�]���f��[�7Ͻ��{o���@�Z���u�m�[CC�=���f����`h�hϳY�Ց+P�+��?I����Ű2�h1pXT,+��Pl9�v�!�c�'���Pֈ��c��Q��מ�qw�S��aj�/ˡ�w��8Wm��<x$�������ÔI'�^�~�Ξ��יq���χ;�:��&��J�zo���|�(�O�V�~�}m�M�����ʅ+~D��L��;<�!�Gu��l�]f�z���z{�L�6�[��O��R�t!"YYY�K���>����h{D��"�R)�\^s7߹��u�9��m2h��M#Ѕm��;C���^�z�����*u����E��m���4��_l�i�8U�6ӵ�Uˉk������D[#$'��莛&�iL��`(��O�ew�n��W �^y�4�sUd�;�o�|z��ʽ�"J�Ƀ|��X8��W�;�5&iW�jkݭ�9����=�:�Bj�_q�����l��1�F�."�B�IMz�s_T�YЛTU�[oD^1����V��4���X&=�i.ϩp�������3��5���m)��ʮ�?�2xf��'� ��[C�R]����՞��"#Dn�=~M�ٞI2n�({-�ó3k?�,�W��a�AC�R:�\�nٸ�}�[D���2x��oEVښ ՝S���r%�< 6�LǾt �-��rM��-1YB����;E�|��;��&�w4դE�/��5�YD�}g��鵐��z&E�r�}���1����K��д}��#��}y/6�����F"lx��(���yMt��׃�[�9�fƦ6��L�t'�tO���J�6�T�� ���-�Z���pڟ�S�'/9��c���9R���0�:2�����w"����#��-[t%݈7��)dP��#�L�<�"}��W^�K��N����wīX0i~ۼ~� �mt ��jGu���Y7��%���f?Rq[]������i�q�=���=�ĹS��KV54br���,�-�W�?�L�Z�~Gw�\��F�����#�i �׭/#��1`���QK�z���4�^y-Kg��q�����3vz8�
7��D	 �|��/|[���g��L�^�cN�#׫���g^��/��V�%�Ⓝ�ά(݂�"�վ
��p
��L��!	*�ǃy2��	c���߾�x+����E�e��;Ť�sNqDȰ"ߔ���0�G�"u��t��k�ӎ�x�j�e�,��R�L�v�~�/�$w�������| �h����t/Tկ2s�F���5|g����g#@��*��p=N�?Gk~��*�Lo��i�����!:Î�x�tIf
v�W3;���G�҃�uݕp�q߲,;�3�����ޭ����()��5K��e����l0�t寛)%�}
��F�Nc�)-������>�<��u�<>������Zդ{Մ7�g&�;q�?�S|��A�r5�	�'[T�EA�/���<�exN��*3�kF>�SL�M5�٪����kye��ɏ�#9���u���߻U;o����?7�G6�v~:��ݰ�n���?Ќ�Wr7���V�C�Ta^
�A�t��Cp�̚��k������jQ��{�ԧ{ޒ�b��kt���Ov��Y�;�6v'�o��Z7Ґ����2���4�k��>���A��t�>!�li�"���"��y��C�\����~4ݑ[U=w�+k�K�7ՙI{��0�/uN1��ŽV�:��9���=���aj,Ӡ���	 �����؀;��{Ey�%�e�U��;	Ǽ=T{�g��ll�Y�ϐv�t�C.KܹЁٮS�Y��d��<r)𶀝� ��*BI����,l�(s4M��]�J��oLn�lG���� ��w�{�ڴ%��F^�]0��������J�~�C�o�fo���~v~�F�ч�z�f��z@`��:9������r�C�s����������t���.�����؅,�����S���̙�s�ԗv��p���.��M��U��o6J�ì�U˜���J3g��4�]���4�[���!�;���E�� *pq�11v�3�����ҥB�/֛��?sd�l�����e�x����6�L^q�$Ȇ���Q��V�ˢ�*Y�H��d (fH���92*}C�w.��W�*����g�X.6{�R3��Ȣb�=��P8C^����C�v�qL�ªh��R)69��U>B�o�����[j ��х~���@����wY��'������_k<�6,��s��V�=� q�"�8����rx����^��|Z�L�4�V^��g�D5���"�x
�0��gI�ρ�(��.����������v������v�?T��䰝yh;\�o+a��9�&Ө�mQ{�˫�OŖ�w^ϻ����2z��+
�=��=�nt5���|E�D�>_Ӳ�,�?�vz^\Kcu"��B=�ɞ�l�v.6�.;��m�H}ŝ�������k;e-���Hs������ő_/�>�%Q��9����R�L-j��*Yt	F�`0|]v�s����i
�eIy�+�[?��\󒞚V�Q�⻱'�)-�0H݊�8o1rn����P�j�v�x�ko�����U"�f;!?.�7��SO	����$ϙ�Q����`sR~'���x�q�/���#�x����ٲ��w����e��윜k�z�d����� G[�n�{�"�5ۙ��7���e��4kҨS~ݠ}�R���c�΋��*������8���?\2�׸���Ιcj�V듥%8���/A������e�af���:�v����o8���]0���[f��^jE�YTo��9��pc��ʾ���b�W32�*�`�6V��NúE��W�[�5�E��3��VB�Bj���F$�$G
�����Jww��KF�����ހ�P߿o<>���׽�u^���sϹ���{b�l`�@����؋��y����k��^f� n�W��-�=p�S5t� \����E���C1R��+�*x�kט�:�}�O ��|^Pz�ܬM�qu��(��;��.Ŭq9�%a��C�m[�;�[q�;����[������M����[���mY��2�<�4!�I̗�o�Ń��r���F�K��=�Lb`L��+�@����j�j�8�0��<�A:���+ڡJ��p|���9��lV����Q u?,���w�̏Ayzf2�����K�9F&T���M�'�wx��Io���G�6h��.	��X3Mz������?�Hñ�~Xc�$�B�m|W;��w�O��xP[^����zW$�9����$K�dX�{2'�s��8�|��>�84���L���Zr�țH�2:t~�ǻxxl2��+ZK^t��P���j�?j���gt��D>me����,SE6w�ЉA��,���uƕ~���X���}+�ߥ�9��o]��+��2+�l��1򶙀�z�O���age"I�"�f�� ?u��B#�G����XWY|p�����P��vH��_g�OFX2����MHS��3?
fȔja��fJƫ�Vm��8gN�4�~a�>����f�i f����KJl淾����?�0�(5��!5F#���']CޭSY��)���ӈb�f�¦̦1�!AQ6�7\�(�=�T�a@���9+	�u�uF�����܇lN4|ڥ���? l7��4YQ�2&8�x��"cQ�'y%<�}\^[Of�i)n�?[��Z�шC���� �R3�i��ڴ�ʏ������eN"P��_�R��R̞l[e��(�PZ1W'Gh��[+��-���s1K<���d��_���I���m<�H5�5T\1L�"�&)TzJ*]H
U�%:��CzM��P��|����z4FƆͨP�x�'���@Dd��JQ�&.�b�h�<��,=��`������T�vE����R-�V:r��ÊL2�_U)��:3�`��,�ZQ�O�~ՑZ����H���*���Bi'q7;1N:�YM�	-%����J���l7���{��X��֙D��Ż#UlA�Lu�F\^���a�UX��ū��5���-�q�9P�������kk��MBY*�3nh���P�ԃ��z�K�Q�FH��JJ/��h!�vn
����R�ψ?�P�p��Ti�M�G�or�_1��-�Ŷ���7����vz��hM+s�����B)k��J��c�q
l��;�f)��R�<n.�W����E���8�E˶�j�	��Iv��:gyPuZ]gMY�pL����,*F��+�A#����j��>fE+�t+0מPζb�~>"h�.cĩfV���|߼�xew0cx��ƪ��E�ז��;�����G=��`�(��^�y~7�{}}S�l.4×ҕ�]�q�����5�Dv���� Z�b?�mt8�T��b�X�����FXw^�.���T����NM*�f4���o�\e���n��(�(8Z��C�~��Tw�J����,|UJ�J��}��g��2�z	"	U���~�CPJ�=7�Íɖ��sC��=� U���\���"�u�Q��FOl���qy��~��Ƶp��{�HG�p��8b��0��Y�oԁ��_�p�&����X�aQc�Ƃ��ǏΧN��W�Z��ȯ���t���>WV>��X���Y��`Ŭ�*s��~އ|��q�8�3٥eTdӖNm�L)��'����m�NX�hr�]7I�����Y���C�}��H�E_���ވ���1�=E2E��	A�0���J��}�-�ePڑq���'�����CM��O���?��&E�LoiD��6a>9[Jw���q�a'�3��.c�y<�<	�����Θ�wa9�����~��yχ��4�藡��g��p٨Q��,LH���*�2FՑ4��]�����5V�l\5�Ͼ
�
�p���	�h=���[c�.J-�����N�|c���x�!�n,�O"o�Ifl�Tm�-�� ^�&!kD�������x�Ȟ{�m}�<�`�5��#G"����b�|ԏ1gW?�$�(������4������&��YHx�S�<<
���Atÿ�2�}��Ⱦ,�S&A�5U������T��-y��ڊq��*��>�> ���!��RϤ�,ݙ�~���N�u,��sD�gt�[|D�۲{�}9�Iu����jֻ�nwµ�BpF"�F��	!YJz��k_��^~ ��6m��Nhr9R�^y�:Oc��b�<�Ps�Bx-<Ur'T���B))B5�V��q�S2���+5�m��-t��C�����ςxn�ܽ�5�b|��Eځ�;)�OB��'� ֊�S��ܸ��I�U<�F@���g�'[[/7Q�Q�3_��w�v"�q�^QЕ�0�'��{^*�T�����c)fV?��*�U���[K��P��띮����;=���^]�7F��� 7�x86hۇ�ǎ�^"�*J���?�F���?�\�eՙ2<[~��x������Ò����� �a �$��2)�0l��E(�/��P���Yfjţ��i ����̻BU�]{�hQ�K�� ��γu��}Ղ�����uƑ�m>y{��ڂ�=iid�v�+ʿ�k�`��Q�j�̚^AQk�N��2m�횕� 1�tQ'~&�U�
j��� ���u|���%V1�$q>5�Z����<N�q۟xZ@B;I��	�
�$���ٜ^}=��5�*Y��@�=Ƕ^`��d�l���C>�-�m��7y	�nR��t=|=�v���۔�7��Ѷ�mL�ɭ��z;�]��N�½����T/7�((4$=��ۭ����d2(O\Hҿ2Ȳ,���=��M�q$+`�/p'�DWk8�D�Y��q�eyU*a���Sp[[[����N�?;o��i*��w��[v����98���v�i��#ބ��}aߒ�7����'ͷ�׸C�^�R�9r�Ql�'�C�zR}�Γ>z�4wm� )b�#�#���RP� ��CwF<͡�Y�W$r�V}R]�T�D���_�b|PH��)h��_�9@0A���ϼ(y�_�,ភ,Y0���{܎9㗝�J(_/�)������x$�7m�z&8�|�� �|/}�酻K��;ٞ���Ӓx�0��u[�5���%�β"���DOx���b��9�H�\�сî�ae�3��3���l���ʔH\B�����}׃r��NsJ��j���O>'$��7�z�G��p璮���nk��/̗��~J�]*���+6���K�B'A�fR��$���������'�8��
��p�<*��S�S�������w��d @xeQP��/���j�M�s�W"�v.���[k�Fμ�R�4h�[�����%`/�pb��b���$0/����(���3c{H0�G/&Y�c����7k���fl{�)��z�vz�1�8��~��<�-��itFKzaj�M���V��hf�A�s���A��\4>�x�|J:qV�
��S��G�$Q�ް�6������s������}>��1�Z���׹�ş!M�������O�k�n��Q0g�*@N��m��y��-}�-�!�vƆz�w�w��&s��ʘ��=�|�+��i�`-��������My��KE� ���$� d�����C�+�ז�Ӎ-�|�l��(��W��:��d]owI.YC��94�D�+OX^kɞy(�S�!�ͷ��G��������U67���Ư:��kխ/ ����Z�T�uG�ۍ�ӫ� r>|h�����P��V>a��+d�+�ҋ�6�fƨ�������v?d��s\��y{_}�E�](�()��4��)����������4������i�ɞ1��n��~*+
�N#义�@T��D"vΊ��@�Y�.�y$����Y�S�����(�Q���*R@�^%�r��s�H^��wb0�"�'����~f#��;k��c�8�,#�]�>���n��E��$7�N�K{��ΐ��r�����˶e�6P�D�Ojon���~x�����?D#�9��[�H:^�`O���%��^K�	npſl�%�0�Gi����&[��`.7�y8��if̙�������>BS�%.7i�gFW-��G�.����-+3�Q�[����@4t�x����o�����Ic��Y5I&o����"vǆ���糿�ܻ�v�6�m������?����v{|��eW�` ����FȬM��g�2�oc:8|\Vy���X��H�T�_L�5�"11l�"���ة��X��t����Qӟ�@��#�ѪbLi�i�g���&.�y�U$�w�:��eP���L�+dј5m�Q�~N���3����2S�O�͏/�M�B��]$GK�.M,g+���m�f��M*�Sb�7+�-wqi�4�U�o�{�G��n��������P���i��h��I��ǎHIheK�.14Q���}>�;_w�2�[�̟�5;c�;�S����m�w`/�'6�:�9H��5sb"�ؓUO%}My�l���35�X�O���i���豈3z�䀅0ywku,j�U��#����ʎ\��懮���7[�^�����������x�/Ǌ�m�B�u��f�Ƅ;���kƱh|�X��]�Z9��+kZ���6��{P��/r)W_אB�3�M]Z!���G�f��� ڒ��h��I�v���"=��NYx|���\i#b*�h��'��2 �n�O[����?5*��֖��*���Z�*��>�^AAӃx���WT.�C���6��2<��m�,4bZ;b���7șϵ\�m-��4Ɋ�ۋ��(�ppY'Jf�ݮm$ߊ�tT����Ѻ'p�1�4�bPa�4��9gK���M�������Ⳕ{ĕZW�J�W�k�"���w���J+c�W������<�"�a�M7�I6TN��z��)~"�����7��X�(&.w'	����"�~j��a��?F��n0�t�|_m��'�23;ݦ*A�~ـ����U�|��Ҋ���+��~)
e���Ee��M~BM��z���5/w���?ol��e�`C���\��6��N_^]��H�:H�;�U�@F��;��%e�=����+Pj��]�D�0��0<�}����d�j*ǅ�^����N�!�F�1�����1��u��A�Ȳ�:�K U��HX\F���5�6�@e�8��4jw��#|�c��d���N���-Tf�,�*�uBT�f���x�\�;[��!�)M�{*|v��j\�:�Km5�ba�jӟ�=}d���;��?|k�O
��I���eY��2i:ZqI��GFF���J���~�ܑKF���9�=���K9�Ǻ_#�os1?�J�x|&j�*���~|�|;��)�H�����V��-	��쪵ǉ.�/�I_"8Dqܿ�0��&ʦC�|;�M�fK�z/�IH4��o�ۓ�?6r&q�^�=ư�������
ֆ��ğ�����9���=hB�H���,��O�����=Ӿ������R��x�cV�����Z��HR�Hy�/�ޑ��+(ڢ�
:�&n���~�oQ�i~�o��j�@O�������n�h�KOu��㕺{d���#�m}��q�Vo9��^��lY�и��{[բ�����K]�#�������������l�+}�t/O<���( ��K_p�o�[��f��)2L4(%BX������8j��S[�a�|/3�Θ42tugm+�߇� N��� �5�=�8�5S�4>±�^�|."�*��=ŞR�2+�[��3�i���A��7�$sK]����N�?�5�n�xc|u��q�g^闕LM����s[��t���s3�W��*�e�wJ)��ha��ʘ������r��S����H�#������z�#<�koI�\�P���h�e���9��L UmS��Yl-~���&�ilq�Б��~}�a"ՙ���� �Ξmi���WǵO՗��Oc�9�q���E��5��*��[R�� ����?����O�#���(�����Y���r�[�%]��r��'��"m��t�ʖ�|�q7��l��u�%�$D^�㛏RTB���$������f��g����tPW����	��yB&æ# �*�L����?S�?������Rl�R��%J���K�}w:&Vm�����<��N����8ߨ�JW���pg�����4S,U�Wn��:�}�����u,��gXWCH�~m<��'�ʹ�Й���Ɣȶް���6Qv7#��i�ǜ^��j5R��`D�^@�5p����2�3m0̈�Y��%�X%�t?�%f��if���1����l��O�ҝ��M1f��=J�S��{�6�n�2
���>�x���7a��ڃC��'�ؗ	�s4�'����,w��f�%�2|�(sT�#7�=+-��E�/&��/*�\��n0i>�%Y�n4֪��]L}��r�\��s�}O{").$�Oڧ��eU}�mʮ6�O�Nߎ$,>(�Cr�6M����[��7	a�ת���\�����25G�Gz��0�>����۱񢺤bL���ӗ��'��^ZW8���:+ZN����lm����	�5R�cɲ�u:Z�~c�w����gZ䰱��cj���:���pҭ�B�_���밓;���Xs܏F#xj�/%q�UZdBǟ�@�J� ��c�@��sV/��'��"��W�Pd����j�n��He�4U���Sꢜ���w�uv��W:kN��>���R�<a�1�nx���#$$�W����S~�zԫ1E�����	*�E��(��v.�#�;Ub�|f�:CZ�y8��i]L���y\eHv(���=�9�x��u�-�B��*:�j(6Dq���̴ۼd�I���,���9�& �)�E�~�0]djj�;RMx1��D��e�'l�Е��;�xF�w��ޣ��m��ڊN��^.�`�ck���#��̻+�Z5��x�l�o<�o-�]Yc3�l��k�m+�p^F��"�T��ɯ��Q:�D�5�^>�M<��M��xn�f�9c���(꧓D�C�V���A�	�5��g5\�/�tb�Ni$���z5gU�~�ܐ��e�m����t�&��y�w(���}n��[d"��}�FH������(����9�mka�ʏ#=�UsPg#xd�R3�ˊk<(���jp��a�<��Ύ%?o&��~D֒�R�ȇ��^���)���>�Y�o�L-�o�{��$���NTf͛v^�Z%Ia��M�ly0+��Ix2A��J�T����i��q-���Q�Ɓ��[O�Ù�`�Y�X��w�f���%՚F���ᡡ� c�Ӥ�:V�￼��X䔎�h�����N5��,�`9AQ<jH�d�>ƛ���5�{�J�R~��.R���S&E�Z%bV�\3�� kW߻s��D͏/�^�}���;u�yd�x����bo2ݠ���V�W���t�/$������5�/{bڝ�Q	̰�O=�c��Yl7�$aV�`P��h;���7f|)�\�y�ta��"�<��P�!�Ea#X]'l*6�2� 7e��b��4��^���Б��b���T�x��CdC�F���%Rvc7I^��k4�I�Hc��L��r*8�=IaѬJt(�<A��&Gl�!ˀ�#]�ᱪiVKGQ.w��F��j	k��}�|Dݣ�r�ݓ���l��~���L�~Y������2eqG��䱿���[�~z��j��j����X�)?r��5�I��\~��1A%�öQ�x쳨����h~Br�Uf�ؼUz��$�i��i0��Ǌ�D� �;7h��i�{��`j��Ng���V_�I~c�RC��/��s%�Y�Şf.������T��=�n�׷��x%��M	Ij=G��3Hb��Z��?��8��=U�
üx����Ӹ���̿�
}�|8��56AY
��K�<�/��V��]l�c(ސ��x������N�^"���.wo-���K��U'%�3���N5������=2�x�\��v�@�a�wT��t��-��`����+W:|���&=������iydy[M�#N��Z+l���%3kVm��? s�E��5�]�[8��p�a$��l�[�7���w��P���.�:�ĵ�"M�Ү#Br_����w�:|��No�"�� )-���U(�/%ѝ�8>M?�vC�>��@���_�Q�t����[��n�㟓�X�m�r*!�ʶ0B��[��H>�y�uvޭX!��!��� S��6ש����B���
�c^�P�Xp��R�}K��w���JW  U�����Gw�P��qg~�q�H�Ȋ�&=���ڝ����nJ���ė��P�����a�4�準��=QUc��T+:�.�3{���d$`3�RX8ۋ�	=�&l��fH��TȢ��y��O��� ���Q`��N��S�Q����i�^�5�w�/�~/7��N`L`Qk���T�����)�����& �ɤ�8�!��Q$a?��R��.��%�g�k}�������V��C�ɭ� ���]�Gf�tb�$`�]~P����]�b��=D���OIK�:�"lش�'K\8�ھ���LѢ�ݎ�g5��Z���`��g
�<�G�bU>�nL��l�fP�ƹ��R�́� ��/�����e��[kw����<�򍫠%��=7ĝ�l���H�b'��[��uڂ@b���7Z��t`Գ+�<K����n�(��Y��k���Ѻa�S�D�v�^���n����Ƣ�H���[49�U�ϊ��L�b�ê2_� +���
�+:��b���uuhKq���rk#h���M)�2$q[�]b�=���徜���4rh�&|a��{lh�]�6"e��M���+3m䅎O:�v��ߧ,��O�e��ȸw5=-�Z���5�u	�d�,�����bO��>2H:B{�&׽���h�xQg���$�~�:��葮���d�����9u��#��dSzŇ�	�-�8>�fe�Mt;�5jJ:�����#�u���Z�R�㧩� �� �f�^A�G�� )Py����4�����x��GH�U@ͭu��;�D�%T�-'�:
%�W�T�<�_��_�hD��;��,���@����Y]��_XN�"�����cf��^O<���&�D�m����ID�V����S�쬐g�P�Ő;RQ�u��5�'�Vb"�S��U�����b�����(O��C�e��<]�|�����.ɼ�V��ռ�F(>�#��X`*ꮱ�	��0���>Mi�g��2�s�(grN(���1��?�"��[��oށ�e^�g`sI�aV�b[)2�zΎm	π5oE����y�w̪�����OU�u N���S1���%�a�뿾.�dM�{֔pel���j�	'h��pN����ޢ��|oYݗw�&.E�Z8I�)į��������[��5{u��,�FR����<�(��H����8e��OT��������d�x�m�{P-Oǈ7�K^���BC���ł�9���)���:d�R9u�ǔ�C���5xIn� h�mD��;r��l�����=�w�ȷP��X&�/����դMx^���T�\��i�E���p.��Ju۫2v	,�ȉnE�mѴ�j�h�[K�g�������[��k������:����K��U�#�w)�c&z��Ǫ$�I���\�Օ*�o��n�ص�(q�"@bͽ�w����_�	���骤M>���ګ�ԟO����:94���Tz��K�>�c���@�P��XCq��h��}Z�=UK�G��S;�,y�3͍&������6;,���}��"����j*|�/�X��Pb�o���\�5Xx�aDc~���X�X�X/���;Z;��.���B���m�;Q�8�\�Ep�����UT�meo4��˫�Oq���A�"�{�~:����k��C�pW��YXq�[�eo0u��.;8ܯ��ϡ[�n��G8�L�e�)��֚?�naee���zK����ȓ�O'm��<�Jg�I{�Z]���{ځ<�u0�G�"M�/�V�Ty���
�ք���9��Sz�R�e�,�-�y�E��r������We~��\�Z�YG��r�D �!�}R��c�s��C�d�rV���Q��:��'E�x�W��!�Ԙ��k�M�'B1G�&>3k�2�#4F��i��=��¥,�aX��������O88�����H�ɐ:E�������N��S�D|g>���+��rیݙ�b�HL#�����:��E��L�/�&�R��>ʼ��M8��2�j�^[�yqF�$�r����#M*��wcL�M?��</RM�@�/c,6snډ�d���x/X��yd�af����S���+:H�(5������ŞR�1��!�u�(�j/yg�����C� ����p�բ�\�.5������(ђI�[�ފ��r��!Y��1�醗l�ɏl���]j~�A����J,�{�W�J�zh��&am�X��ݙ���o���2s)��+4��97Rݧ��9�.�Η��ܢq�ɵ��<��d������TX�I�D��˷��>�D�R�����b��ˍQH���ƩY	r����,0&v�\�
KNH_T��T�2&g�:rj�;��d�G!*s^�uа=�4�2�%��O�g2߰���T�j��q��Frf�CU���D�G�pzS���׻���""��[��,�J��蟅�Ћ}X�z�H�`�(�j�hy��R�<��KIۓ��&�7���ٕ�3r�]��n=F����H�YW
A&$�B��5C�����b]6�����=#��߼���ﲳ��Fk(���:=�L^��x&u��A)�z�hT�J�#�XE�����`?���z������rr�cz��͘���7Ό��y?��u��P��c�Zſ�%/�zg�D�3��.+��0b:�<�������D&P���tZI6�����]p��$?>^H-c�l�[S�M$�`j2��j���%A�4Ӂ��7�})�۪��ϟ_���[�����<���,,�B*��`w*%J�Dx�6V]�I'�X!}�F��9�`�4�H:W�W�I)�'��f���LA�As��I��溻�/�y�?������Xn�N����3������P��/�-u�(�{t��{Պ�C9{
L�.��-X)j���')�� �x ��C�,G7�5��� X��ؒ����!W"W<��P ��r6M�/�ëټ7��h�Q���}�μ�wFᝬ�vt��0�� i��a}�|BM7��O��O�ioo4d���I����WW�	^+��Dk0%����hWp����g���r��Yw�gKo����G5�/�t�~$s/�����<|3�1���0�D K6�����Z����-�R����x`{�:��	CUC-��',�N;9Q�mEq�]�R��[��m(���2���M�\<�&���q��Y����fj{q_�h��{i8�f� p}��[�n>o��o� h>��&?�������O[�+gq�������)�T�����+h��⡿�ͬ��(�uk9��������,|Y��(�h�	�����9�>
������C-t�MЬm*��]1-�%���f;==��p�%f{c������)j���c)��Ei�w6��滔!�d3%R�l7�Ή�-0��v�_�����;w�z�����8kz�Ii^VY �b��G�Ũq�N�d��#O+}���[��n!btܗI��
�&h���4�\�4�Sn��I�1{�VL}#{<��i���䣶{\���
��Q��n��ߚ�:����"b�;E}�	5!}�K|W�Yg3W�Km�I����͐G/�W�d��WE
�O6��&$���V|- ��X�����O����j����;M~4������qHC�o���7����
K_�~�O�X����#��y����N��ȹ�B���O�8�3r���o}	s��N��%��YҼM�72�Լ�'��w0�U�'&���=����?�9"��Hk[�@f��|�_C�T%�÷ǟ��e�Y���
U~�\0B�]�m�����mNL��������38�~���vr��c1��ƃA�ԝ��/�oI�ѐ7�8<*��\#�{of�L$�=���������:���׆����Ί��*H(�#ض��m�!�\a����9J���5
�����Im�DJ�/lQ ��U�R˜��<������	(; �6�t�q.�9�
CZ?8�=tp��+��_�&)������0/��?�4��x��&g.�FY�׶7>O6�U�߼�I���X�������1��_�]�r\ƾ�^��'�\�q9^W�?���7�QI��u�{O�Kw�di���|�S�s���g�o9 M������=���� )��-Q�v齠|������=#
�op���-��F'Չ4��)�r��w��*HS�L����PK   JrX�@M��  2�  /   images/a3f7833e-13f8-4e96-ad38-aa22696f9742.png�y8�o�7|[�H�"di����Ki��-ɾe�)E�%d/bb�%����c�Qvb�c�����<���{�<|GG�q���������u^t����� A�ʵ+���h��w�'<L��{��q� =%���׊� (gP��%M��߽�����I�f�rͨ�����6G�0.��3��g_P8v��l�����+��8���O�':�ٳL#��/Kc_��\�U���wu~�4�@{\�{c�
��=j<]����˯�U;vj܃H�d�k��ghe���,�UJ������/84��!���Ϳ�˂���xiSSӊUL�G�����4q��w�ou4����7�:V���So������!u�ݻa�^�n��I�Oed��A���h�5�P`��[uG6������7بݠя�Ү����d�2��W~mcy��ˣ�a}�%DE����"+���G�'vmu�<Ƞ!���O:�G�'r����P[�<f��ׁ�'����Ms�V��iE0�?G��!��|�P7O&+]�:���h�K|DC�.��Z�,#z|{��#���u�E�O��Ĵ�H��WU�+����n�/Xo�pgC�J�8K$���b��m��
Y61X��e�_�ɫM���J�����S�>\؄=�~�޽ӏG���͉��D�t"!񕄮,+��E���h?�����"�w�ޚ�x�#�b�H��h�u ����u�K,�%��c�4�_Uuכ��Hӌ,o�f���:�T�[�����b�1~�G�/�ǟ>}b�7�e�w�Q�j�F�wO�x�ެ�_����u��d}�gL)�,XPY�R�K���<�h�)O�-��c����S$j��pHV�0'��"��}d�m��n6M���^�N�v�poi�c��m���\���Ϻ��u���Kh�{�\Y��B�����֥�~�q������K�y{���l9׶�?~|ȥ����(��얰�����}b�}����X<<��zm卑��;ʉj���S�I�@�3,X,���̳{I��O�un���Ȫ�EG�<'XK΅��Tr��j��f�}���6T3l�\��I}k��~Z@y��.����;S�PM}@;߯� �lH�IvBؖV,���1x�y�FR��ԁ�t�A<~x���.k`�̱��l�P�]k���+S��e��ꎿ�?�Bl3%a���/����=�H�i��O,H��V��z`����%�� `��`�%>V�ANZ���i�51��.=4Uvv�::E����?FXS���ZX����99] Z�OI�=w�-��}y�����ə��Hq���bȡ�<Y��>�U���*<��q�Ϯ9���o5aެ����8�@�x]�K+ 	��%#�`����iy��y�B�o��R���'�X�y��d���$���v�Tݛ?ћ��=�xps��g���ʐ�w�1�\Q�呣w*H��j��g��d\���9���t7�����J�/���{���L�G[��bL���3��27��x�v�}G룆�\�/p���Ő1������ N�#���f� ���Y#�$� �˒t�S�s��LX:���,�(�5��OHl�c�u��;��������GF�y��G;�]��x�bf�}�bځ����g%Lnn��s��ߨH<�@p<��%^���΀������^�~L��v�U���y566�M�	����G���qX�� P�j'�9�v��6�W���Ivy%��,7����aڟK�l��X�(H�Y*��L��1�S���CP�8D<}�`��|k����A+ڴ���T��Փ�6Ω�b��>�Lק�����V�K{�̐����RܫнHc��K]]�xtJ��;�,���4p���#K�+�����W�O��|1k=Ǚ(�Z+�f�x��)))�XHĆ�a�w���t�^s񈏒J[����0Jl���\��{+�\��Y�[A�+��8Ų�J6ES�j`sK�ðڗ/_L����v�`��OgɊ�c�i�s����[���ߘ�##�����RZ�X�����c����������Ą4�~���2�{qq�E
6YYJL��Hl��`L�pp���w�ڦ�J��ϱ8�SM�5^ͮ�G٣�.��u��0�X(����ٴ>��:�Y��)���EH�����>k3uh�UYx�a��I*^�=����(š��������ރ�>>>�
��Պg�E�Y� .ZI�N��\B�}�p'ҿVMIb���j�]�!��9+ǵcb!K~y0��b���:��o���fQ�nn7펲�\�e��c�l������������3a�+���s�%e�9,j�ֱD{{�'{��5Үē$���<K�#�;�eH�vwrr��_�Ԕ�⯽.�F5eU�(���H=v����e�Lo%���k�����/8�<�%�����[�s8�WR^m#���R4T��&u�	�����xx�
OW.Wlt���'o���󣛾k��}�n����>�m�Ԑ�4�&�k	�Hi��*2�_���1I�s��D:�L�N6�Yc���5VRW8���Ȫ�������N�sl^ ��Fc&������z�q���g��	��4nw�$���sMiU2:��z8)��$��D���;����y�Z�zlr��mps1��
j�Y���#���4�Y۾.e�{D詁�I�Z���H��GH�������ĢJ�e~�)��c-����)��7攔F..F�� ���$�Of_7=_5�,� �ߢ�r��iI�W/�������n �R_/^�7������o�8���<�.���RF��W>	�>�x�=�(_����E��O��M�pMs��/s����N��0�1�vDBJ*�._�5/�|���ي/�U�I^��HkOsKKCM͕��{��{O��/w*$nR��d�ͦ	���A�n"���t�$��>OTߺ�5'�[�lI����&b[L�F�A�<�ҧO����K����%�ɱ z6[��8�y�Q�V��`�f1raK4ɏJ�8�DwQ����Uz_�Dvk�Dh�.s�Hd��|^�Hx����(��!*��/_:����GP�ٷ��b[���!B6�E!&''�E]�v��}� ��I�DD�ڎ�S��?FGGp�t�te>nС�q� ?�8g�&�k4c��p��#��F,��EN��;=HW�>q��������K�����Q���Z�X��]�e;ƌ�y�z6��y��Zx1	L�)��j�>�����ז8�npkgV��	,�m���Z����I�"`�TD2!6=@�A(��v�n��ZZ�O^p"�\U\�P���@��[}��[\�|¨��e�u���=3�Т��XZ?�0�����[e�f�ܮ5�,�y{��ي �Vvs`����k:&ff;��F I�����LD������?~�uf�b���?��֦]�����w�`������Z�N�S�V�v��y�wA�Ǒ� W}o��H�L�PA�Qcc�<V�|�`,�}��y?]�b(
�W����N�مL���略E��ظV���n` ��Պ��5e��;�Ji�s��4Q������������O�����B<:�+Hao����@���hg���z�d����A�#�@�N]	��� �.�9�<t,���(��I��F������A�Lٙ���#��n��x�~G������/��s056���r>��2�;d��K�SE����s��CYIR�S�wOq�YAv�j��ާ^��D�4�)rs�Y���L���R�i�o�ؘ�lB���VK�*���(5�;,gb�v����$���떺�H�}n�{gL�v�Jp��PR��!g�O2s����` .}��!؄�4S��i��*X�!�=s_�=��W���� >����ֺt��_K�%��h���~�5\Ʒ=�ЀΩ��l��脄ȴ��9�!��3tVx�~q���;���C�Fک���{������ i�cɝՂDjȡ+(�5�]i � g"��K���nF�>Ȭ���Xk^tČ�8'Ѿ{c�c��ĜhF�`��7	w�ݿI�{.�"�R����A`ҶAG����8��g���&���5I%;V2���[�291��S���ɬ/��Zeڷ����kڕ�8�E��)�J!�H���zʫ�|�`�m/��U&���[������La��U�օ�>�i��8Aߞ�<�(�l�׋��I���BCB�So��B�Q�&I~�7��}Z���1�Pj?V�p��V�* {���`�n:�c"��s��n=����&1��~Z23�[6,L�X@���JFFF� *H��V���@#/^�x�3�(�<F��9sR�gy���p�O3�s�hR0l��Ҥ����뢓���]~�ctf0�xק�555��V�c/��N�홲�&2� +��g�{x�<��s)�v5�U��^�{o[���ii.���V��i� �q7��"�AU��t�A��� [�G!	���'�z߿�l$~}�2����?{�[{V�W!���I�(�"�� /���<��d�������V�}�����t�~2ٍ������ܜ_|��w%���{��D�(�K|ͦ���4m#��ͪG��|��C�B~���Ƞ�=u���)xy�N�u�Kf��p����f�V��oF$U�G
�(hj��BV�Y�W.Vԁ�l�#S���&cC��Q��oe8�x��*�������y��I###��El��	�勥7��׎�w��S�`bb����8�Է�\��l��"�Z�	����ݓ_�|@Hu���j�(~�~z��I��)|~��@�q�~�MzUr�>�-;TG	J�=��o�&��$%
�#W�����7sss�b�]���݁�� ���fJ*6`j``��t�i!�R�M%����]�yy�l"�������nڧ��m&~�њ���Z��-�����-4�Ikv�����;(�����z�(3U��6���A�@Dn�3/K5���߹���Ձ��\9S+,���	C�,�=ǽ�}�r�Vtpy$1lJ �EA�*!ː�W��,5$R���S���z�
�[F��������z�x֓�FTގ��$/e��^�w�����̒qA���&F~��`�iy�gs��5�l5��M����.�R��C�I�	la��(dD�[uݗ?�{�J�+�)��ӯ���Ӗq�
ٿ"�����ˣc�y��5$�����ﳂOl���;�7��K��]���Z��L���S�����ח�F�EC�m�f���C
���񊊊SO\k?���p,a�n��W����p}��{�+(��Ⱦ�r}��!�rm��I�]�!e\;�4�*��aC]����ÄӤu����ULMMzlY�Qq�фn�����`�ɳ�2+}�s������--��q�=8FG���D�m,�E�.,6��ܖ���2�)���'�9�k캡��o]�܇Ji�	j��s�*��D��{���ߟ_<�{θy;�gǲd�.d�R�\��nƍO�>7GuA�y��V��b���4������������i��)A�f�����bוui0�D3�)�:O���V�c������˯v���S^���R��	�޽;
�W����xuy�nC�D��|+{=�p�X���9GG�Y
��жbٔ�/?I�Goۘe�h������x�H]~�})e �J�Fl�W]�_�WG�Z�|/�[�4i��N\�(�Dǫ7�(����!`���a���ȕ��C&�35��r�H�Xb�:��!�V.�>�f��h�O��F�|b�Oj(�mZ�2�J,���'��K}�Q	D�	����-��Ve�������أ��٨檱H���e�<��˵���Q��������G�
 �\z���v&�v0M+W�L�۠�t�5��=~v/9����x�ƍ3+s��Nx�ʜ1�6c�2���׻�Y-`�P=6%`W�3 ���w_���a�u��zwj7���������I)�>zZ]F���硍c�~t�W�.6a1���ዓY ׃7Z~8�}9�ĵ�8O��j<�TE9�g��X��t]���MIV����}Kŋ?���S��l�]�+��/˫tؙ�׃,O(�ȸ��;�4�|@����6¥�WI�VV��9B���H�[<
����m�E�������[�����<��l٪έX�2��M�'n|��8Z�2�;0he�ڝ�)�g��PI�(e0X�b	|�XXy��ץ'��
��3ÂZ�d������)�P� ��>�-=�^�\L�]�/\yk�}kk����'��b_afSU���Uc��w���Y��Y���SK��Rd�����L�h�s׃�� ��3�,�U].�]-Ԧ�!���8�Y�%l�Ĺ����e(��6���1��l�B�dB�I�CE��`�W��b��N<����p��Tk2�,��{=6�$o�g��������}�C����y�����APra���w��YM�U����[��U�},Rr���9�@��ZldL�2Bz͵�����Nא�}6Yq����e�/� -\wJn/�������h��ĕ$)��|Refb��ా<�lW�9�T����`��b'x��}elLu^DvH�4��HՓ�����B]Y�����ò�~��?�z����O�o�d�'�d��(�R"q��AxG�d�#e����U.��i�r�j�_D����,!Sh�6cB�����Ǯ��+4ؓ"���kVsIY 0��}�g��=T�6�7�&��ey�@c��t�*2�����d�0����P�>�ȶ�)�Wa����S{S�,��_��a�?X�Ļ�����O�M�k㊑�\�yf3A�I���仱:$d���W2km�4�U?����c
7I�,����
���F�X~M�,�=��{M�ϯ.��_�W�b.<٘	�&n���j�X@O�88^�K�J����o��'���av��\A.��s1�6��'�s��Qe�jO��K23ղ�+Io5���Hhoui��W�%���j��m)Q��+�~��]3��F�-�����vo���E��mo��T^�0����R_s�U�.�̘���.j{4���9�J�$�O��U=j��|���=����&&��Ls�qzo]������ole�Z�ck��/g�����8�g�H՘�W��E�X���G9\*$���Mb�o;���g5!?����x@�(�Ñ	����L<���4���p���ㄡ���j������g�p���t������#=��g������e?w#��Ka�y�5'���WN��4w��32PL;�֫n���|ã���KҴz�0e�E�IH��ڠqa�^�P�$K�}-���^;q Qm�ʧ4�G&����p�ƽ{�~�	�����Ync��Zs2��c���LoK=M�M�<��k��ﱚ�L���tL�s�S=���Ǖ0��G�����C���0���u��j�዆~��.J
�Z��ү~��QƧ��,�w>�P�+�]��H~cm�u�W���݂�S��zK����*a�ONu�����ui������'�e6^N+���z��d#~���1��^�}nf`v�~݉�{��i�ML�Q�L��ӗ]��Jr��}pP�Dֶ�׭.E1BP̾�:�Cvə���`��w�j�t���n~�����%��i��dTOx��:�V�k���XE�3f�W�U�Xm�I�uNZ�޽�C���V�	��6R�F�ʂ�V�0?� �+ԠQ5e!#�sڠ܀�3�4un����S��@�a��-�w��Q4Bu6��˧!\wD�{�T'̾)F��~�P�ǖ�j��)��)��dg�5�
�+��<SP�g���尟J���%^Z�c������5_'bo,��@#CW��|��'1ʌ������@H5��p��4rxF�^$H��T^S���D��ҥ��W&�M�a���[\��]55%.w�ܗ��,?�أ�؞�u�v��v�wi`�'��1��&)*0i�ʳ�t���	������x������ܧ��-lm�D���^�<t'�S�0��q�J��l"�С��!٧�@�B��i��^um���|^԰t&���n:�߿���Ʋ���q���܌ׇWן��a��b��Ģ����>NY�_i����J8BG�����O�r�ј�/�i,�jxX�쵅�޾L`��PXn���K,^_�|~��xD�-[c���Ox�)����+�>�Ś�^���]�"^���}��5�� �Y߾�U����� V�jh==~�[�DCNK;-�H�&�C�?W�g�:�Ww�+�~]�%k�XEKll�����LK��]ŉ�a��Yd��_��O�JH���:%��'p��մ�@r%�v}¥��P)"U�&�|�/��Q���ø�:�������ZQe�����ӑf����訇�랏��n!�[����Լ���GZ��?̦����' ��
�Y��νZ�s+7k	 ��K(���b��&d���V3�N_<�Y2c�4cKe�kv�b9ܟn�y����sÍ�Do��ʖ¬
]���Ҭ#��XR�n�������iu��'k��k��������]��P*~�s��<��T�9a�i����w���T2lZY�}��Gqs�,4sL��P���#�<7�KO�� \\��Kcm�������D���j�:��^?�5T���~*�1N��Mş|]�\����m�B�">[׏~+tP�~10�����ݫ�p|x��G�y��N9�i��ӵ.88=L�X}Z���\e�M욵�Ϋ�) ��$$�����{ս�H�%ֿ<����ңA�V:*��|)y��$��c������y�.��ERT�{|�(�����j�~����L�܏?�7�c����*k�|�~|����E֬,|�uFr]Ϸ\�マ���WO ��9s#f�lb�?H�����n��9���A�p��E�����ʩ����@<�'�o�W�M�RT�F&^z��N�T��~��O�K!x�~L�M]��x঳φ���~��w_�j������
9K�k���0'�3*�Q��`��p9It�@Q$7\`G�h�1mM$�r5q�'s˜�A�zp�9�M�b�]i�r]��R�Q��;���}�aF�UK=Kӷ��LgaQW�C)�򓳔A��`J�|=Z7�!��d=`��Um!(��v�<[%+��t�f�w�Na����WeE�E}'�Y�W}ks�&�J6=T?���+�U%�[b��EC_|�'\���r��< ��T\�j�!�\�"QOEjrl�bߣ�RT������I ��QG�ˎ� �H�.�u>��/����1�Y:�x<����3��\v��r��4��"/̷�@�Kʟ��璴}�[ꪌ'��.^�ny�>6λ��}���SQ���:��TG�.��I���=������d��K��7�J&���ȕ�c�����N�+���BϾ��a�T�GZo��n��
��e�܇�����>XP1�Th�WB�+S3�
-=F��F���<�}Ƌ<�8d��$�;�� \�}��Tԃ��3�L�WX�F�߹۸��j&tvv�|��^�Ƶ2��t�@r����g�V6����,X[oMvhՈ��W���{V��H�N�>��M��n�vT�2�H��z�A�x�AhO���?�&�-�ŧv0˃k��s oB�ƭ�Y[�gk�%w������f�12��	-:	�1	o���ݡ��Tb���� ����b<������a2�� rk`q���Z ����a�T�éOQ�)��x񚝍M�I�h�F���<�q�fϧ6n	I{��%�ߊ������ɂ#��^3W?��=Aw4û��FC'��5�ܤ(S�����m�2Dz��u�?�)�e�zx|`���g�#���$i}%/�
�WI]r��t̾M��	��N!�s/����񉉹��&b����>cs��4O�63L���gq�3��~�<;$
wF��6o@���{]���'r�����}CR���/��Y

sR9��KV�d�z����"�p�P�HDK��'Y��H�ƭ�b4������s����[J�)�9M�D�?y�c���,��7�t|�:v��O$�����b|���n�gu`��Q	��b��4Z9�f!�@s�Ҋh�X��Z�q/c���xo,��K]L����*��~�w�����T@�.Ү�-�du%#֣�q�F�o�6����H����-����sL8B5!�$��93�9u!K%ޅ��!����ϯ����?�ʱ����[��'��#Ezm�;7���vp}�Ϡc�y�'f�9V���p�ḫ�7�*=�lNm(mi�Q����6Oi�z��O.�m�iT�*[ed��1�Y��w�p��}2�ߒz�Ӊ��P�a��}�Hz���@�8`kkR�}���/B����M�'#+JΒ	%LAe!^����샴ӑ@�Ŧ���W�9�?��b�J�p��_�R�����p݆�ۨ��̓�(~�Z���B7�>ĥ�0���]:��n�{����ٱ���I��E�?��>z���lg��L9r$��͊�d��Vq�&�f�K��*Aa.�2�2��
���[r�������>����٨�E��)����0�ơ�ڧ�auڵ�9+z��C{QT^a\<<rY��D;�y;60$�X�*���!b�F���M�P-W��U�����>��o��%$�~��[̘vK�ya�=A��?<I�=�5��E�j���Ɯ�G�Y����w0�����䢋������x�����f�БdIS�3A+@��Rڴ^�<�`N�k�8t��v"o�WK��aA�c�,��Τ��~E�����z��j��! ����������1�|4�SD5]�v���m!�n���{��*�P������?J�0�]FFF���{�������S0��G��o�_��贲�r@Wz@�;�c�<a�G��
/XP�66Ff�Ú~�-��5��vsJ�L�X��;���T|G�UĮ/mm|�
�:؜x��G9��g2��y�~8���ҫ�E<5��
|ܕ�)M�'�6I[0"��N�E�T7h����oq��u�~H��;�}�X��gx�$���j�h5%.,�8#P-/BB������J����[�,⑀��;Ԑ�3d�<��c�Ζ�}E*EvQK|��*¬=�Zj�k�=�Yj5�����[��U�/I�%���M3���wI��q�ԅ5��=}�~~@bF&+�'�l#$e*�^�]dɞ�G���H� �;�$�@�x�
����ٚ�S�2ngc�wY��Y	���q�9M�uV\k�]���l�t�h�1�-b��I� ��O�e�ӟa�nO�z�Ɠ_�M���Sҕ�!�r�#��4����q�%����%��j��T�ii�M��	��'�%$�U�N�L�O�|5椫����E��ˋ$;�.�D|������M���ˏ����1Qݳid�Ш[�{�d�u:�Q%
��\�*dfM���1�z��ߕM?�"8~�!�����>�9���80�����lUy�ؘc���oi�Qڧ����B Aj޺�� �<_�a���?�^L�Tl�\���Y����(�K��)I$Kï��_[)	X���`�ّ߿�*���m��}��C���w�b=��૮�1Jp����*��Cg+� �T�P�l��>.ƃ��%�.����]���7I��a�����ؿ��37}7�;���
H�|�����z�}S���2��8���W��c��洹44B,U��_�^����� P����b����[�	'�z� c��x
��H,�V��R���5���+��wQ� 9�U����}`�P9���Z�i�p�	g&�8^��)h�'B#�ԋ�Z�+�x�� D���*T֗!�H�%A�ǥMO'D�Ơ8���z�q}�M�3>tR��d���vV�V��j�(d}�e�d�Z��=�|�f|ֆ�A���{~�}�����@l�C��R�G�s�i�0j�_U��H��d�x����
v5N�..�9  ]A�mC>����l ����ۤ�Z�ѕ��ڡ�|5�x�x�s/}*��7CaiL�x̛_H;`�u���Z��3����P�h�������/�<�5v�v�����dL ]��
h���+Ԯ�1��fE���� fm����]evw�}4�zoү��*a"TO�x�xW��l�7MS0.��f�ڀ�z��c¢�̱�g�Z%��*��ޠ+I�DbbːrDzs�r�&�P���!�����5\�v2���q�p-���	!'CQl\��q����IUWi������v��3[G���fe��9u�MD�e�g����g���80�_���tP�MOO�O���]�;N�&��XS}f����\��f��4�v�J��rr�P\J)w��nDw��+��G��&<���zW�<d)�|��)��+髧ix��f�S?W����� ��j�����jp���h5�"o/{�Je/��4��;���>X!p`��h7�®c���D+�>��U��5 [��=���7C��h<����E[SS����=n����h��Y�v�;B����ǿW3�[��6&mװ"��#�۾R�Cx��zo�8���!�lY?}��^�^hr^^�����R����
?U�Μd�h5�/q�/��n�r �F�2q"�1�?��cW@ +7˽C�ob�mgdH��w�P��6/��#�D�|�ؕۤ?�\�M��h��ߍ���R(��s2L}��^}��-�q��Q.�g�bR�Sy���� ���~:��^r4�ۍ��+5~Ǐi�թ�VN����/~��j��	���/���4g����"|�,����ڴ8���n�guq�?6�����Pl���"��+Q�I�~�^��A�E�6ϕ�5��o7�z��e��l�ף:��S}�:R5%�!���u-�z����N1!0�h`r8����?5^Q�����ԣ\������J�z��xC�0� E��߿3��%C�@vӺu8�����T�˾��k�BnվT!�0n)?��9��K���zHX_��a;����*��۽{�U��"�{����Y���^~�bS�
r/Y��Պ�:���*�?B����N��b����t�Wy�
R<��}��� ���5tt���Y;�I��tl�T�/˭R�|�˱�:X�IQ}�t��d�ӧ�z�4����&)c��J����[K��b�Ch�����~��H_�)�\vc�D.�BIs��XP�K�Y���3ͥ6z�u�H���|uuY	����9|��h���
r33�Z��%��v�*]<0o@L�͚nmC����j�4���F���*�I���f	��ق?����8��{�ȏ����Cn��{C��Y�Ə9�v�y;E<F�O` �6�ƍH&�÷��w��AnW�e�nP�|ޟbZ����b
QNg���Jئvn���_JѨv(��*�(�. ��5��ojL��pa>��~1�q��ߋ�����G$tAB�J�h�Gp�F��&�~�<�7}w|/��Z�f&�e� ��2�)20V��iOs�o��wpJ�*�;�����R=�(���&�ݓ,���t~w"��*[��%�vZQQ��h[(oe0J��dTV��������G����u[�fꗪ���w�O:����0a���v,���KC4
s�@� C�)��Q�N'Vo�V&5�G���w���|�������\;Z�@u��k��Mcu͟P[����S������pᇿm_�}�!���iȣ�kZ��w�E���Mc���J���q�}�f�
��������Jf��ع�8��^��A�����9iq{+�4��F����l�K��� Uޯ]79��Ḣ�3�Y|(+ �w��6�f��u''~���t�/�ݲ����_ׂ��Pr~��~d�V4�B��l ]���ֆ��D5n|*˖��9�}���j��p#��饉�������'�L(g���.�0��~::�,@�Wep�?W%��D@�7VB�?@��S*��7n	�ӎ*ۓ�5Ҝ�t�X��������2�H��2B_�Y��)�SC�ɱ��?����eڻW��iP`ŗX�,�I\OѸ5��}�֯��P��e˻n���$�H�ʳ"�#~J�t�1�> ,9��F�t�����(�s!�Wh�U�[�F+�~9((:�#:..��Ai+���8�^ �js��_.)
�P�Ɖ9��ޛ�Zb���v1��K��>�]#{��0� �/w�RMAnɺ���%j[|�y��N�����Z}�m(�����m@AȌ��?�h.���u k�����A��S���n�{��#蝻5�=�1���[��E�T���qT��!��v�g6�� ?�y�'���ύ�o��ǝ�n5�P׉T$��X��y�L��v>nyy����;�TMA��������`���Ӧ1���No=�3�"�˺�W�@.��G߿}�w��//o�q���ڙHUL[	6>�܁�>b ���Wm�D�a3$X͍#s E���K7�Y�����Ի���U���^_�8�y��]^O�Wk��NA[XX����}�`R3
��=�N�:�[��&�����ML�����ѝ	����b/�g���>4[ �};2�(�,���?b�+�P���
��Ǿ�xG@$�C�v|�&11LЬ{��3sGU�?�A8�9(I궃|�_�亜����/o��HzpwjH��Έ�I�g�-��>8�P�d��D��[b{���~_"��C��@�:'k�����`rٖ;��G����B��K�Ɉ2��w�옝��1�;<	�N�H���y+TԶ�u۟8x����95T�g��1 O�'��T��ظV�䏺+O�>�&�>���Y�s��~��w����G�>~�� �3;ʹ�y��X�_a4���&�
�\�1�shn�|��I���
F�AT��Rxa1�������y��P]�%�����/�\��rJrH�H���=�����ii�<\i�A�-xGP�&��"��훦���)d�ó=���n�!�����!��[�֍�.-5�p��[��U��d�F�wF݇��UTUl;�B�BPh4�6��C��׆뀫|��ԙ7��w�&���a�6��&�$')c1 �"�m}TQ�#��PO8ؓ������ u������u<�~]A,�w7�q(V�	�G&�_���C��%��A�'�*bJu��6�B~BX欼����]ʬ���]�D������[���&��jz�N���;�6R��Z��*e�n���/��ǵ�|W��*��Y뵴ҥn����.[�Wb;|7��T���t^�ء:���5��r�~nt�-uP�I�ۯ�菞x�M.Q_�s���t5N��E�V�h�{@�%�V�n��$u[^K[����Mo�%C�B�F��t%�3/.h����J��R�8����|�8�����J����3CR�a�ҝ�Y0��_�D���t[(k�J�����L�Ȼ(�l���w�U��<k [�S��]�4ӛ��b��,��t���/8i����S?��ڳi��&+�c��|`3�|�ji���.��v��<����j��	����ͣXMC��7��6�X(�B�wf9j�R10a��!�缵]��&��!yZ��j�zl>t2�s�X��H:��O!8�6:�%���P% S�^�L�?qq�\���v_v�df��F�pI�`ie/��ΘA�n��Sa�%f��5�zz��}.���W��|?J#f����9�|����(1Ӄ��V�Q��y���+��V�C:�ĭqî\�pj��p���2�t@2�8���$q.��8^]^�hX�ѧ��W�F�����]�-�θ�k����z����Y��4�~C����)��ު�-\�G�F��r�AȦW@���[�G̈́����X�8Χѷ%�4��d��m�p	���=!���^�^�,�oE(X��_V7	���2-9v*�����{�o'�㨾�¹�[Ӽ�a�e;��?�}������
<���:��>��ޯ�:,�8�D� ��b��u»;�b��W,�;u?״Y^�wB.Nnu�Q���l^�ZA�33mҹ���C�k��ZA���֝��xȷ�{�߃�����_���!q�Ǯһ�'ۘt5���S���]�� �4|	�j�*� �>õ����8?h����Be�b��Vp��eg��Y��_��3�R929T*�:��	�c)db�$C�T��:\����R�g�r�m�/ɋ�0�,	S���g�K����aÊ2�������*?)֪B���;C�$w��@x	��x��%�R̋W�J��P��H�v�{]����>�?v���͵%R~�56K�������o��W�K矐�Wg� e�t��m��Ʌz��������]:����x*�;L~�LiU�Q���C���6�c�L�o����6���� ���#>_8��}�Y��ȡ��ag���T~%,U��Qz�E��`�xT?��,�-�v��Y�x�MZ��5��T�	�M��+@��y�]6���Ҿ��[1�6���ݽX���x�:,G�.��x ��P�Sn�9����Yt�>�`�yăW���|XO���.�����o��g�b�1��,wm��y�|�C_�Xj,�ʋ'K�۴-����l��񭝫xJ����t��v"�g;��G���DE����Z�0K����"���� A�=��_�zWT���o�u`�jC~?��_��=����{�߃���� �MK��i"w�ʝ����ɷԺS���N���8�0mzs˥י�q(�n䙂Τ�8D�Z�6ð�"�Nn�����'�rv�y��-5n��XQ6Oʸ�x�WM��<Z����
�[ا�໾\�x���(d�3{=��k�k(�s��&�2�Ѥ��Q�!Lk����o����`(���C��KW��ޏ>.�Z��X���W(��~3��;�]f��ϲ�?�`���	ʚ���>������`�Z=xD�4YN�+UK���{S��=ie(���n֕}O��3�幑��5��|�:�2�����F�J=��g���a�(��~fU�I$ ��]��r|�e�t�()�o�d��e�|m���ú��s�m�rNi�����fR���WH��b�����Bf��(�Y��C�[�z�N�}~�%�.Rj��G��6A�RY�Ae�N��¥� .�S�M�什~�?pa��&�7�I�̥;ϻ�l��d���]��/vc�K'�3W��~7	CJO^8�[�ላ(%U�z-7�Z�Q���9^Ct�����Y�:�Js%���܌O�\��v�s����Åǩ�/V���Syq���d<�yN��[�_OfЪ�*s���vU������(�µ[��S��~E�!~�ɒt�����:^�2A�gbL\W�VZw}�������3������]
��7&`sO�Q"E��o	��Fh�yO�m��k ��D�J�����<�+��rK�����+���$3�M�Q��w۶l�K6 c�H,��+9gk�Q1��v�(�M4d�᯷�p�>'���P��Z�i;��&;7�.W�wc��b�C�$3C���|��	�v�(Cw��h������i�Z=�ɝ(��L�l4��T��h�]�+p�$W<z<�*$�:2�/P^~&/��
n�/Z�0<\��/��?˼1ͬ������ J�T)ɀMX���bʩaB�@�����H���hY�E�J	�
�EW�x�FJV��m�~8��h�=�1�J=*=u��R��p��\.N���._��[���IPS9G�{��O��h��q}�0P����V;U������{�5���� 8��6�� EA��X(J��� ҋt$��Rt����P�I*����W�% - ��I��s������ˋd��S�羟��vg����+Y�����F=��!^t�ߖ3��A��S3~�FFد65~,r�)�O��O	1Đ��q%+�U~���G��ǻ&i)��²,�+rX\�{���oTX�\~U~g�M�3�lM���r�At�{�7{��wDȄA���G��GђS~�S���]���mq;�]H9�A�8v	f9^I�1�WO^RZ�<�bs��\���\��?e���� ��:b�S�YB���wO�k�◉=�)0���n�K�Q��S��̉�J"��YI��C-S��6�Q��D��z'���Y�������,6*EN@m�g"����N�os�N1�]w��yY��օ��ܯ{1�a`YR��d!�]�R����	�~�V�ｇd-���_uLl��+1��A�x?P���E7�kװe������g����w�k]�A^���)˻a]�����h�fo�Ж}���&����h���W��-eT�rN��0+ߟ9^#��1r���vCo�B�]���T���&����:�f���K��ߨ�����K�~2G��>�"w\�~��㕡���ܨ���G�$�t�7?��g#%r/��+-G1j�=��f1��B7��E���#�Eϴv�&_ύ���XHm;�/T�čs_s>�1 MkTt�l�-��y�lta�\��\ ��q28�1Ja^��V���l��c-��1AoB��9�9��{���I ��.��q/�ιj3��Fol�|�)�y.B���P�է��.!p��xSc�ZĘ�¯�g0k�J�����n����[�Sw��<�Tk��f�W��y;"l#'���h �W���$�J��nƐb�S;��H��DSBɯ�_��C!J+˞�W��:�E����	���*r:���<k�༦&�w�y���Ǯ+�!�O�%�m��U��k4)�D�.�1
�b��3��ϵ�'}Zλ��I��c�&?�t%M���bD�3�2�}%{2��ʰjsi��y��S��eՊ�Q-�<����Q���a�X����>�O�]���..V��� �������m�A�9߅��,f�}Km\%ѵL��'�"���z1bw��ظ�둟n�uO��d�!	�7�[���۴3��������핪�ɫ�T�=�ZQ�G�kU�a�غ�ۃ�לB�J�l������:�M�JsH������<!��5$ka�<vc}�k}iBU��U���:��Q: �O��);%�k���a^ZŲ�'ri���}g��=M:�d|���~��	�G��q%���!�N�m���e�4ks}�LVRS��jֵ�F�x%zfﰖw�p��}�Ő8�!x�8z9�C���)��H���<,�N5_���}�U���Z�{f�1_��Y=��Kм�(�Ŝ�؏���"!��~_��9�`ۃ�;���z>�K�J�v���~�UFEԅ�Y+v��Z�e�X�;����4��$�/�ߝ��1���`{���E���Ыv��~���&Ԍ�4*m�?�pBz)����
M�*$�!���0����/-H�tۛߋ3j����ƞ�Zۦ�5���ݧa������?x߆��ٿ7"Y#�t�WZ �TFX��������;\f��mB�i��ά�}eg�}1�?�L�>��P{x��n7��M�#K:5f�qB��m����xr"� &8{g�L��i�e���{�u@0宁���jGƐD���֧'T��'ϴ�J�?�=�{9LJ�jԀ�a�T�> ��g�C�L�WN�;^ñ0��J���L��ĸU&�W�K�Q�ta�
)�Z�s�C��3[�G{�9�9#R�6lZ���~��s��ٵ��c��{�T���W9C8����ɛ��z���bo�(I$c h�,��YmS .�90�d����9>g��j�k�3�N�^�N������ʩ;���٣&m�F��t�G���j�6���'���n�U�G���q���'rșLǶ��"��O���;la�j�b��F4��An��Թ��p8�poq���e`����}�Op��*q#�?�6���wP6ZOJN�Yj`��L�V��H��6�����˞8v|y٬�>'��p��ed�i����f�P��Y0�:��¸⎠�3�����ϗ=����J:�
��a��w���eh�������aʲv)e�3Y�Nt�]y'�ʩK�\�rىB�tC=�4r:O_hUY�)�xJ(pE&Pj��8�U�z'b0��V �C����p��%��~@��l�Q�]1�o|u�1�?��j{>(�@�D����e������|��ayT����/z���U����zc�L�L����F]<�;X���xt��a������"3]y"|*-��%Cr����'p0�H��MkiP��%А���"���y���\ۊ���U�/�.��|=���5��J�CS��j���q�]�q�k>m��%i�<L~^�ȼ����/��L��w�'z4��r21@�lMV�w����#s�}����:R3�D���*�ڵ��ڱm��N�1�on��~��.Rv7��)�;�[<���r��D�	�+s%ش�_�&r2"��H j��d��\���^"y���Q�8�b���F�ԟ��[�y���˾=\8R(��AvM!MU
���K#�5��K���9YiE함�tf�}�K��,�F�@���O�Y
�R���T	�4�Ijs�	�u~�)<i[k�^\���P�������n�2���a���.
Q��V�Z�Yk^gč�M����C���N���p[]y7���}N�_���������b[-��\qK}��2Q����s�]���<����yW�[�es ��i7�GM��i��@�'��(O_�CN�n���K��T�Y<�����}��]Ŷ�<�=�&�R�"w�4�,�c��wN>9���40+��S��WY�m���٧V�5?�ޢ�0��.��₞+Gc��Y���V���*s[ɥӬ����X�&�^�1�J ,<}@�Y����П��&>�u^�5�G�zo�<�]8ϩV^�4���`^�aEP7������mR�����M��������[OM74�V�eq�q�w��3PI�[���l�~k�m��p��+v��͸�ɹS����������ͬ�A���@��n/?��=O��ݣ��A����K�����Xk�F��/�I�=V9���.���p/��y���7.�)Ё��u8�3��Jf`��������_����C$��1T�3/����0�\C� j��u�}���p�	>�w(�"}��&'f-��H�`�*�\�_�|�?񽁒�W�y�d��*&6��?�!��#�d��f��έ�h�Տ��\�����=�ִ��1��Y�X��C&F�U��&�>�/���x�	\z�o���U֑��u�'���O2��^�yo*�W�FP{<mz�n��͘2&Þ������������}�{y�?�{�n?�u����2���x�zU̿oV/��(�#W@������Z.���k�xPp���&ɸ�ԡ��`b`�~��Z\�f��G�9_�����ư³�R&�*��iκE�6��JY�D�\J/�-���o�)W�Ǉ�~㱳F(_�?S�8.qi�a���É/�K�=�6�x0����m=��}�|�T���(&<��N$8�/�"��{�!�7�BI�
��_m�h�N�s�0����J��ª��*$x#I��2��~�T��s������n������2�g�,�œ�I�C�b�TVK	�b���fL��A��/�s�Od"}A��A.W�9�)=l���_9@��P�8���^s��C~�sF)��ԽC���ϧKg��5��<=yɰ�����9E����[�%Uo�︜���Nt�?�v�<'�m����+J��웤!�|{ƌ+z=�\R�`�=�mʫy���}]�rȑ�����F� ����ض&��q��GXg�y���
���N�0p����t��9�X��E������'�9tx<P�}1*�7���S���]uٹ��4H�p�����]�N�Jr��Gm�D��&�J�bn|�@�c�ɾ=������Ơ3f���%�!f�E�%�i����xM ��z7�f�k������R-�
{��XP�*��dnO8Y�$B���}��?E0����f�"N���&�?���XX}�[3L���v.�k`�lND^�nL�B�V��-�:������u-Ruو�f �J,1ї�ced`�������{6�,ّ�%��P>�P�G���;�b׾���&�@#Ha���(�.L�xzۛg|"�fn3G��=���h��| ��V����%3E˹�I�$'a23��;�w���󂣖ɥri,��}�T�ln���J�[�BY׵�=�+�ϷD���y�в�5��G]Gy��X�ȱ�����w���E�vW����Զ�
??�����}@P��=��C�e���]&Et ���]��an�ݓ�Aq��:c.r"C���b��P��w�d��٢���.g�]�RV�+�
�{�黍g��6�8��7�j�D��-N�c�+��9��>q�2�:�ߝ�7A��Y�|7��s�^����˵�l�����IY�@�.� {��Kr�������`�{�+F��M�{�>��'}�+�Pàn`�f`�h�
(����77=��$���'\���*�D�����M�ۡ�u��G�H��(͌���r���LL�rHa��o�w�l�;ڦ����mj��v��^�k�	=��=&�b�IS��S��h��~�ș��J�?���mH�Wu�U��~���gp3h/�����a?6�Fk牳����{Z鈳i0 �����H�9����-�n�u���7��`���R4�ٍvQ4ٻԲ�Nw<!T�_o�P9Հk;���l0���۵<>�71�R��P�� [��BD���ͳ[-�u��7�)���Ώ6	�	�S�2�W��2��o~Uk�ho=V��?Fd�0ݥ�;_���� l�Wa�vzX!��\�����"�A��n�̤�:�-�s`��/'��'��\N��'pJX(����w�t�;�'X���M�,���*.�1=iUn~n�Z��?)X}a�|s+��i|}�1[,Ho	�
����-������"QR��Ak�W��a�s�{1�e+�)�p�g�mC�[C}Axt��$8K��V2p�Y�������a6���0��}�9�V��t)?#rl��ն�V����Qe�T� ��G� �_9͘�M��g�Wٶ$ήR��Е�LJ�Z&�l��	\���SW%���= p���~8߆�aaPس��4N̴��g�@���h$ȡ'w��8Ə.<;jwT�BK��|a[��H	׌dK��J|�c�ů�Ծ��+i��u����I��Z�e`H \_x�4|�k^���.>b�S��-����|��W�Ƒ��0���LÝ,�J��5C���u�\n��s�T����=��h4��Z�Y���Ч��}<쳪�ֶ7W0#����?�ڟz�b&�,���&�ڗ/_�
��<P:5�%��i�O��?�(��lK��ox
�/��t)S��@�U4mj���ާ�P`�8�Z����g���ÿ������+�^�Y�\ؘ7��Qf��"c��=���O����v���]a����N�~]���n�l^�Bk��Pdd
�#���qU�99��M�#.��̯�|�z��+�}���R���D��&^�Ŗ�9LU���L��X��5u��|� �����H�AW��"�ԩS�)Ĺ9�USl����_�i�P�iFGG'U� (k����gt�RR�J�EQ�mmmZ�V�\`�Z�lyg`�l����7��yF~��d������ΘĮ�������b]jj`����v�l�_o��]YU�gddt��_/>t\�����']`��Q���M�=�L��oD4_���p'W�} �W����m1^E�B?�����_�F6��c/�2�/KKg�U�<�[\��6��Hn�@��s�\r~})�w)ʯ�L�]���������ݵ��x�l��
�ui��)��K�o��T��^xD�M%���r��602/u���*@�� �[ifv>>>Q���L6}�c���}�h�N��R4>榩8sKG~5�9\ Bq�,�2���шZޚ+�!��f�5p��G�W��^��Z��e����]�=Z���oB�=����Q�S,�F�7-����G�.p����Iex�I�;,���@{"�NM�	�Ƈ�L�f������d�$vga�XwZ���i5����gCCC�ee�sz-��1f$&%��/�9�h:���(9ݏ���!ʤۮ �0��kdA���������T��,&RN���lf�+%��Б�2�����mu�[+P���b�_�>�e�f�{m�c�pb�J���Jt���[��/A��T�­+�=v�T2��o�`�\Y7�� �v��@�Sݏ�����,�[s��9}�a܎��>%��q��C-�kR���yӶ��X��J�Dm �<�	�e�����[Ri�ߣ�KyF5y~����E"�g�R%y�'�o�A��Y`���� �0���۲���������<+�Sݪ�uK��I(�KKA���l���*��ќ�2�� H��C��!'. �z}�S)����h�v6�5kWf�۳�g��� 5�
zB��7�O.҈�k��<��T�^�s����O]5#h��|���>4]'
�4	�iA���9 p���h�����q�'\��Û,����}��X�,ɡ:�,/��F��Gi��Zp��]Se"���Y�)]�ņ5���>w{��p��w$�D��ޜhn���G���`�f�f?%_���۰]1�����?�r˩?Vɛ���lW�;/��5X�A:�r�L��˨��Jk��|��ڍo�5�%�s̖2�R�n���'cM]��*�B��[�H�wzJ���͔@9,�>Q��ͨf�3�z�a��u��w%�I~W���Sc�6��~8h����� ��`�*/��t����=f ���c��M�~�}������x�����һQ�n<����[O�L�n�	�ǒ�?���vU�4g�b��K�)�\2��ތR�$3w����=>�D=��J�D���iM�-�iv7C�%�fU�e���v��?�.���-��������҅.�hw�s�:c@uE�E��RGGF<k^W�Ǹ�`�� //�B�5�!���۪��H���P��pS��gо���Q(�83�[E$/)+F'_ߍ��7n�஌�*����w~��� ��p���)B���j��R�+��k�.% L�<�Q),eN]�uD��-�kR�Vc8`h2�?r�.��&�0�9��D!EQ����t���5��"ŏ�Y����%�������M���;��	H؜�'l�P������l%n�	g�:$�=�Sd �kg���B�Tm<r*M D�y,�Y#����>ϥ���%�0��
�ݥg�Y�������sa2j�J��U.�@�ֹ�cz�s�S������m<z�T�ұ�3��u������-�E��h�Oc
�j��X?�1�|�.�� ��$v��ڙw��(	vHT/}��,6��Ʉ"}��-ݚ�ҪP�W���lF(�x\ڋ o�{��k�$��-��5uxX�{T��o}��L)�]A��Y���;G�G��(�Ӈ�w�?4�����͆w�^:m1j��������K-�Εԍjo��F�f���t@���F��?gW7^�E�s��D8(�=:U��[I�}���G"��#@�ν+n�CP���μ�z~�jW����ڭ��=S�s������gE]�6��q�����T�������쮈�Zl�qqI_��;�)�J�Վ�������2C� ����݉�����	�{���M*)�*y�M�[?�)��[��E@-�7wŨ��5�:�]���%�QC�V����ms��� e
e���Q�;~|c��O�y�9o:b�A7�'9�A@�6a��S *�ox4�<�'��mʾT;v����5܉��7��פ����ռ3695�5>>.���J"�o�n��qRq#{��V�q��*u�N��Z�XDH׬�u���+	x3�ت|�L~�`������/'U�EsH%�VW�����@/��I�J;8��~�Ў0x�-b| ��:Ǯ���	@�*ǔ��H�$n�j��{Fyi�3KjQY)��ȏ?n.s�D�Me��������ڝ-�i��%Ƚ�������Q�8
�IB�72x�+ng}5��:3���cW�-V�W����ȋ�yȴ/6%� �ِ?9�<��ߨhۻ�hX����6�|Z�R�2nW������0��i%D����O��L&��s���������.�Cp���WZ�О�2��h�ll�n|+��i��E�'�Y�Y5��\T^�m�zK���*��n�B����;�&���p�G�f�
��ᨆ�S�#�f]�M=�{��O��k��4�,^TTL��ai��*cr�ߕO�X�eɊ[�C*�n6"���l<v�a�v��c����~o�]��Լ
�zp�ޡ��~g,3C�����R=�7��
��k>Ԭ����Oi�h�F׬R��3y��_�n�Ta?�5f #��L	��Y��GCFF�
����	���F��bT�z�^�� 
�BJˡB�*紂�.�F\��UJ]�?�`��[���`��GO�
�\Qjj<��9�}e���f ��G�`�B���\}��l�\TTt<.'_0�jv�{Cv삙��a�Fnt����Z�;�i����U�B��\���VӅ�KQ	Pפb�.�a��gv���l��:���zi&�'��]��4�t��m�܁�\�
��{��;����\��sEQ(g����K��{�(!?��И}V ��0�Z;0s&�j5�������v{��+�@�{�W�䝕@�h���opD/��I�wft: ]7�kdǍ�W��-!�)�.�&�wĔ�G�ݜ� @���jݡ}Sl����ޛJ�S�6xr� 8B]u�P���������i`�ܩ_]9/��:�t(!j��9/Be�/�6g::�������5/�+b.]W�,��T�?pojLRf�Ϻ/${걺�$����=�ӡy�� ?A��e��z��W�ה��8!,d�]�A��,u�2R>yM���#��P���0HL��K�Ml��S���wܱѭ;��ԩ4x���f�-yH�r�3�n����+=m9w�x?@�JGgPP~���n蟥>w�-�+&yQ<��$����s�z�_�PfX�z2�N\�kg�1�WD��Eyq�T��!7Y��`��
��ܣ����
¯i5�<lJ�G|�UH��	�&*�n�(� j��ChK5�_�5]����VWB��Q�ą��/���o�[�A�����%ƩD!;3ڡ���E_�Wb�tn`�]��Ǐ�>�###�8;+�.Ι��������·[� �j��S�=!�U@���_�f������V+��8��j}Q;��T�cP��)י]�S�	+��,�@� 7&; *�
ei���9v�
���j꣔g�;���ęJ�H�R�\Ks�1�ąM`�Dhʽ)+� ��F&�;lƿ�|�o�
%ˎM�ߧ|���t����W��w���3�jˢ�g~F��<;�5����|�� :,^�7�~\���F�5��p�&���.{���f�3�a�-Qqs+
�H�d��5�j��
�>��`c��m�+o_�0	ʨ��ni�K/S�?sE ����:7UͺƳjj����y1)���V�,��Y��٨�RRR{�ϨE�{PAz�?�<��P���D�X�#�(��q��;QMI���v�� �X�ڂv��� -��j��w�-�җ?���K����rF�sY���_i��n�\�ڷ���u7�w?��I��[�~���t��1���݅�v�V;��P�?�_�ԹT����M&�(�E,�"y��w��E��U6�� 4�ȱk�{0k8Q����V#�����WεE�5Z��W3R��ڛ��_�^�
7n:u�/ �R>2"lj|k��쨤h���b� ؜QSb?�v5 ��>��;&����x�~A;ِ	�S�~4�}�C���@�sG;��э�PcGǝ���35�]-����ӻg��я��a�;��{����ƚ7�<� �#��m��fo��tDTTvEE�PHbé�����h�C�e��掑���;���2��ўZX�2�7����ٳ@�NL�q�6��rU5���c]x�~�2�'���l�b��镋ўk9�M<2-5�bMr��e���Jƛ�>������˒���y�J����9O�Y��ȞW`��!��Q����Z��_��;�ʁ4/�S5L����{�1mȷu�8��]�"�S


/���%����>��m?G��5�}o��Js�H�SƮ���:���?��ey��̦�.0~���I\�����ɩ�����78b����hk+����F"��*��cV���HRRa���?���%�� ���t��h���$�:��H�������Z$9wWJ/��\{�G�+j	v�d�� ���*g�غv鞿j��*�h����V�@�8Ea*ٳ�gu��?6�n�O�O�;::�f�e��w7��6b
�Y-��G���C��	��v����x��K�n��UU�vɯoN$����kG��~� A� �Ĕ1;[[�;��;�T��ʤn��'����ʺr�F�X׫:���x���tΟd�������.��~�{l��l�=��$�����ҿ]I�U���&�̉~��V�9���^������`R1uS\�����x����fff�Ǯ���L���"18y��4"��.M������%���ˁ����)f�X_�ߪ���9PZR���<?����[���YS�4
o���;;?���q�M�8�̧׋T�y$;8:�?;̫���P��h�ԥ5�F������|��w{?��������՚)9�\������Lܕ���EFR��/��z�鎂"v�H�����z{{��mm'��2.;ű�D?���TSS�a��ID�FNrh���0��_&�3�)�����9�[T��\~�~e�A�������ճ�6�<�X\�� ��������~��+++*�^�S����k����b���]����[���dx{{g����`�����/_ڧ��E��ʿ211�E���}�c������"��! m��;����&��I�Y\��ot\eP�����\Gg�+��x�G;x06�aø������Zz&_�&V�Ԩ���H�;��S�H������1���%�����]�Ȉ岴����h��c��ס�\���Y��㳓!�Ԩ1�����f�/jd��>��N pE�NqswX�O���.LMoz�|,v$�	m�A��"v ��YI�P薔�f֨��M��I�!�
���Y�m}�"'�$���������ynq���ak�Q�_���p��WLe�����hhh4�s�u�UL�NPH����O�P��ˠ6v���FS� �;������I
�K�`���x���mY�hSɃj7m��7o�\��R<��;���NO�`�LC��
����e _�D��S��h�-��Q�y�NIRA!�}��*RSS���j��aB|��3g�8��9!*?�1�C����F`��Й �9�:9P���|�PҠ���.�2�� z���O���p&�u	�o��k�������������
�-�@�ONN�Y����cgg�+b��5�u�1��\���������;��AR�	�A���ZZZ��`�F0>���5%9�Bw�a0�\�⨧בI��_������`��~� ���x�,�XzJ��";�\jw�P���!z��ӕ�(��"oaA�X�򢉟��'ii4��8=Y��f>{���&sy�%KG{����>د-�~��TQK8�2ޟ�VqE�.�m�&t�(�߳5����_U�$��` �%��Ɋ�8A�5t���S����z��������;0��a��f��pC��a��� ��l5�F�>�3/�� ��,A�D?��S�W� �����H8V��<��� ��CI�U�������YM	mO�'����ǐi������[��qq,�9�۟�Ė��e�(��k�7<����Q�,g���|�+Ն�����{����ERJJ�_d<���秅@S�r�T��1�2�&45��&4A^���i��qE|���#P"/_��*++��b___T�$7�`���6-��� ��(b�Q+�JK�, �c�F��cK���2����;r�K��F��B�_��'6_���� R����I�UU�����EA�ei�ȭ|4����Y�봋���tZr� P�M�<�&�r.l~&�"���)���&&�v�/��Y��3�
���_�x߿�1=�0!M	��������|�xh]�Ǳ�.�x�v�'qtO?mJ�-�|rH����9�RuQ��)�!�+PM=�����1���h�kl��4��uS� ��#�\\���q�c�y:�Yԡv9����B����e��`0��JO�|�Q�����+���k H��O�@�h5܄�+��Ç0�?��NHK���jS9Li��)�Oq��Y���w�q|a���p��R�{sNP�i����� �g|���:�CE�\Md�g��]���0{Q���V��)�s�da���vU���u'� �XF=?5%�����+�侥�A� ��MZ����
:k�=�i���!t���H�R

��5qo<� a|��4 &n�@$J��w�Ґ7莰ބ&����ؒ��� \�;���6�6����X���ل������ƺ���'$$X��j'�=�#k�_���*y0�cZ�ӧO�����D��uv�~q*�Y�-ѡ��$J��sss�-���;�yM�Q2�BM�FFF�>���q��b��u�-���n	xp;(�M榦�� ����~��3!���.>,�ԧNA��b��=��W�X��'< ȫ-����a�!�
�
�"���Է�xyy_��l���䢣���> � @귾�Zd_��/x�˩�j����vJJqN����mG���~b�X}��R{o��ϸHuk㧮���r��B&�i�����(�4:#���=ҺR������~'����3l��b1H l`�b��c�^��s�:Н¾���ﻎ��TF��^��Q����m͚r@�@����<��h�eē����.����*�~�aB@A��EM�4����p��*9ɀ���D�Sp�83�A�r�Y:v�lo\�s.�ڲ��7.���Z�V��IP�='�6!*�ӕ���M��*s@8�W%@��Y������\d)�5d=��jVu���ŋK+�����\�j�(B��^__�z�uĊ��|��['}B�����w:`���
��Q �\��L a_�-�*��]bR�ޤ�� ݀Y���QO04^�V�z����XZ�������K������P��O#�?��%4%�~�ɼ� \㯱NɣBw
��~��v����X���m����F��m���;�Φq����� ��K�ݤ���oV
.�z�-%�߯^�� �.J�ռ߮OVi�n5��j\��J�,���&�ӪDB���}�	�d�U;!~�3�x�E�#q�kk���� {�}��fT� Tt�N����g�DMZ�ݞW��ߋ��M�6�]��
�P���њ�[��6`��K�ѿEoU�QŔ�]�c(�b�iaT������{[EM��iS���^�����U0�ʗ�Z �`;�N?�����^��ɓ�j=�su� lTy�ed��靉p��ē���e���L�Nk�DW�ŷ�j&�Љ�3�)Obo���N%{�F|������I$��N�WC����-ܐ��)��^0�o���MP]�6�s�hR��4��-j �`��4���;FO�N�n�3����(�3��D���53�wjJ���۫*�AhAEɚK��-Pb���Ф��"�������!@DjHLLL\���~I*�(IK�@b �D���iy��^�]:���A�T~UUUN򷻥&;f��+D�u1����qj��/	������"ٳU�@�N�T�vV W���PB����<�;�Trg�����?�3/]���qF���o_�|9I�� Ǟ��@_6-iJ���Mk��;��L"�5��(Oh��m��\9;� �.@�hKx<�Uմ�V\��j����<t�P���\��Gy��#��}kft�+'�������
D-+v���uc�9(�s�,O߇���2����f=G���.0&
��� �����_gń�%�=��D�^�<CήM��t�h)Խ\����G��<H<��������"k0�#��T�޼݁�����x`�̼��E��#=Ӓ����k�Y�6 �@-��ń�j�T�	vw��8%ew�ƹ�dPO���N������K�Ɛ)�mN@�UH`x�����zx�^)���4G_��X1%Ya�	��ۜ��C�L�R�a.7��)�T�����P����u�D*,�|QUQQa��	um�X�?��C�n�z
���z-e����H��P����T��({�z�MW.<��}i�2@�3�-�3c�Ы �Z�"�}��y:/����#��ʊ
���t��мV����������ԫ�F�[�	>=m�R�7�����sL!z�{k`J)�T��p��X �R�����������;���`s�a�E�^�+�]䕽������L����1)g����I���k�j��Ih@'E.�ZZ�Z�+��x���1�.)]9�.���?�LRڨ�OP�HyG�+�w�~C��@ *Gh0��
d{2	�Y�HV���t�N��V�|�^A֪��K��G&����W�̀��|�v��{����44rY7�a(x߉q�~���O�)�?�T2I�����.{TH�S�x����[[�&��XGʯUg<��)b�� *şj�.*�4a?Z��/���ʙ*�������������m�
dP�����p��y>"2�!�ѱ��r�l i�~��y`HEU��6�������]�}��vJp8�������#��3� ZЦMD�&1�NY����d�~k�Q��t�v���U��k!�A��x���nB*rR��xd��
���s"��V��Տp�f�>����D�u�� ������J����67�}�U�e��)gbV�l��(�M/ٖ66g#��C� ��c���x���n���9���ꛌ�>�q��G�vvh/+I$c.����

�}�:C��0;� �n�	��?��m��SKM���y� �[W�׳ �zu&�PX��r���`N"�詩��..��zZဏ$i덅n���ɨx�(Z��x2E�s֚I^�h�&�I;#����ј�Ud/M����͍��)�E�^�F���K�GKS�r.`wKY���Q�z�h{��?ۛ�@&��줜Q�ܖ��D+¯���fg�
�}*SRZ� �"1M	<wK���~v�6�7u������џ}U���СL@_U�iv�/<���j�|Dp�-j<]�>s {(
6@e��)R(�

�*��@�����B���j�,0ߡ��H`y������)(�v\||�:|���R�� �R �6�=ڴ9�y�����'$X�]�j5�	���јN��2]��Ӫ�s*pp=���8
i��H z⛣�iK���?���hV������<8i*
���Ot��ݤ/�	�m��d�FT�7�|#�ٙ�@�`v��Y9�	Í=��oۻrѢ&O�h	\���tM]������NHS�42-9Y��ԅO��C��D"N�єf	K@ ��T��0l�����mq�ͥJ�t�A��	TolG+(���q�`��p�Q��=.	���&� ^.��vJi-��@�����u՜n�K���ъ���J���c��U��q������c���Rv���?��ݸd�M�\Ԣ��vŦ9�⊻�[d2.>��f�׮M��F�ܧ�n津���鎶��v	�s.�*(�*�oo|~Ɔ�	�5�-�U�I�z$M-�<)1 ��W)2VѴn]Yh��4��������u�pÿ�h���	����n��'�	E�)-��{i��m��<9�]�->ƭM�0�@]�򰵷?�Xw7��A�����wT^����A�L@��j�٢��y��6X���{Y�8;���2h9�����	P־>���;�w#T
�"�%遦��xW�S��x6�?�{w2�l�w4�V����H�=JBE����3��S$���S���כ�ii:r�4�*e�&bC��u�"v��U�Ϛ���]coӢ���q�ߝ�)c9p�+:\�?z�YC���z� J��e߼����|��0�v�3)�O�PO#����[Z&p��P�SR�kH��?L�h=�Z�ftr�"�������V��:m"���x<W�a���n�QO�ɹ"/��+)�
j�����PC�s�zfN����f��x&u)��<��	%vo)�������H<�
]��q���ǿq���&Q��l R)���������\��Y��K��)�A(A�}��Q�����ed����B��=��a�� �K�P�m���!j��=���#��_+C�!oB�����If�٠��6֐[UUU]W������T67��m����$��߄�E�qvIU�MO��0h��b�@͡/���:����w0	[�4����~Aql)u��\��_�
hh�H������P�9;kV�b2b�i�%I�m%K�([U1��쫮V����^8�hB�l3�E=��!0���K��A�4�����D!����c�T#���kk;D�Bm:�*g����Q�VI�<U`�ڔnӺ�d+;�aN.��Ɔi�~g���l�'�f�;U"��{�G�);3�i�������E5�.@Y�ZF�!����+>�Ua���\!�����.�t���n�:�#w�`�U[�T�5�J�
���y�0��
y����w���#n��׷�sS���(C��Wa�k
w,��x"Q0C$R������e}��a��t�U��a��0)���r3A=���p� ���������3%���ǽ��r �����
�Hs�f�����j���{V��F��&{}��1+pG�%���)j���i�f󈊛������hhf�'�î(���Kç��j͟�'����D|ᬋu���JjJp,�/Z2�#6�u|��u�>� ����3!B|�s�R���o
���:�4� �ՋG�-*�����ҩ�ɵM�P�Vx�E��=�ǖ5::��������tZGzד�_���f�ץ?\����KEc�3���>���t���~?�@]�gG�% {�ڄL(G�����ͩ�/S�>J��B�P?�(����g����>���*����H ��K5�eZH.TRCI<��?� es�6�T�h=x��O=-`���P�$;���"�ZGh& Vq>:krr�3����4�5%�`��漦�r����E����r%�gX_��Bo>�	�[����utosD ��=r�E�����8��l���O05M�UK�!���� )IH������@\}�Dгo���W�Sk�5DP��̅�&[�8�X������f?�< �x�~�ኴt��t� ��/g����:�䰣�s�O�$��h���BB�fP��� a��s���>�7����9��Ik�J���A�9��Ki0:gڞ� ��)�C�����u�c���/����`�w,ꯆ�އ��a���8|�.C��\{�ਛR|#�Ro�fNP�MZ�?��FYk\�:����p,�=�ʹx����|ؘ��qK�Ԉr�bŮ�(���'���u�o]b_����g�� �8�%�/r0Q+�p���i�����غY�?��\�L���a��������Y�{���o�kE�����.؈��rZ�!#�DV^^��0�$a�7�[���F�d�$ K�;$N:B�R�Vοn���PK   � ~X`$} [ /   images/a8bb870d-02b9-45f0-bd60-404fdaa8f6ff.png켉;��?\_ϣzR�'B�OE"b,-�����f�v��Rc�Z�P#$��R�l��3�c�Ⱦ������{����}_׹|���9���������u��;v�Ӿ
7ܱco	�{77��'���������O��X�y���[�;D>��wV;�0�Bk�D�ۡ1V^�;0�YG7g�����Yw/�D���;��І_�����D����,.����? ��?v�@ў=r���>?Ot�8���g�8�Ko��ve{��;��M��g�d��&kܖD<Йpo����k,ѧގH����@5F�G|�X��9�@�j`S.�'��[��ؿ���\�m�݇m�h��Jx۵9w���{�D�c���W��%\[����vn}����ma��������Ƿ}>�cN{��!������	�#�{��.��26��������.��qDSx�v���61H�~���/ڈ���V��|~
t�Kk���!Q츨(��?q6��k>�4�r�K)�TnG� ���*�E�Op�@�]��\�;/˘a�y3D}?��J�������%�����ٌ�<�U�Rb�pT��f�%�\��$S��J�d<�T%6��#AZ���ǻC�zs��0���?Y����z����c�*�9���ޟ(8B}�Uv��K�!���W�DzS�ڿ�¹QFn���\-�-|�&L���X^�M֫�-�d=꼒��t�?�>,�����3�ah�1 Qf��qːY�����)J�	B|U��"����;h�5횇�p���7x��-���"ǵ0�Mø��3j�3��$���6RɟVS ���Y�|䟇e��&m���>.�E�{�.�Hd�Z`����)�E��w��4	����ۦ	h��;���b(��?���3�nԛijiY�7���[�f���ʢ[�M��-o`+��]�S���ḇ)�˨4�`s��ϐ�5��i=ΩX��\��0�żӸ����Kpx��J�e�ztW�J��erC})�� ��s�>��+Ȭ�?'�a_wu޿fg��0�*�{2�as����@ۈ̥/���pK��~p-j��uۖYo*�%H�Ab$rp|�,���6�FX�0��y=�M4n�G�'�s�_�e����>���x�d�k�������f��$�D�����=��_;#�z���c��$w�����O[�&�V�
��?�ݾ��|t���A��U���à�Ϫ^&��A��uص���qX"����
+u&��SJ�V4S8(�}�")�+��i���k�<j�~-�=w����1#��5�E[�ws<7:)e�wmt�U�#g��r�1�jB�{	*C��/Z�X�����V���E�i��Z.���E�pa�L�PS��<���w��C�Q�S޹��G���)!�*u�nˁ7,�o�n���b�:u�J�����f��A��J��'.f����O�-�g��8B��$�PI�7u���;����z�>{V����K|��Zy>A5c�
/g����1�Z)6T��|�/*��,����MD�8֒��9��++�����4�`z�Mک��e}����ќ��CYI���
�Z���ŤTe0-�FY�=8����E�A�]c�uc��^�/#��F�R��kqbi7�jԯW��U1m�/̏��bh�u-m��y���W>-�2�߇	M�H7ڈ�2{N����b%�뜈�M<�S$��r�Ot��e���K2ǯ*�|�í��������'��k�������:��a1�����J�����������&�#�&W�J�(�bUOx�J<v����.��rcqC#ĉ_�E��f|��%�h0L뻸�3a}��a�k��M���<^���~(���`'���"k�	=`��5�����^�o�EjB m��h*��ɡ�{_��'x������R���f�����Zm��f�4i�U^��AT]��!���Q�UZ/E����ÁD�J+��նܰʶL�%H~�;�g��ƢGF�L?�����ť}����ōϦ��?ʱ�c�����d���^������k�i���IL��@�dh27N(��ԿaUJcmm�O��y�w=,0OL�G
��;~|�*��Kc4��M�7n��`�c\�����g���Q���I��Jg|f���v��h���)�՚���mr�)N5ڤ0�e�X}���{Xm��_�ƺ�"��%�#ǚ�a:��$m��ŗa8�$����N�B�z`���|
��q�~���A����ӻ=jić�Q}{s��6[�
o�J�$���j}�~��P�p54�!�3���A���F}�©��S��C���q��9]�OPY�v��r�Y�0�gD�0��gLm*+�`����pS�lp�����I�2�rP	~!�̕ߔE�<F	n�g��a
L�)ݽn��}����B+	e�h�s �u�L�j���n�t<,�M6S������-�2_��+@�p4�Lʾx��^����p�U���q��ҁ�}!��Ya�� �Q� ��ʪ�S�oC������������l��Okx����m����V��S}<A�mH�\���E�ֿ-j0D�:�̼Lڸxh������e�T����Zl�\7�I��n~�b77�N5i?[�SlD���6��$�pJ)�>x�ܰ6�:�v��!�	��J�"fz)QÿbJ��@��N[��niI�jZ�N`!=>��#o-(�W��\�:Β���	�9�qyӒ-t��4��v4p+��a�7/yF�0�#�j�;#�@�_2���q�B�J�Be�p��?4��j��n*�����3_����j���*�~��v���7���m5�i�!�P�V������P7����;~�M~�2=W�q6RkP��*��Z�>r�&Xryk5,�6�qJ�ϖuԎD�z�K��򥹇�+|�XP������HY_�(�X�ԭC�Λ���B0�������c��f�M,;RP����vQ儅�&Z aa���7��F�r�=�Qu;�HN����a���6��2�\��,Iq�5ăj\���n�OPa��)_Ɏ^P?���Iл�CS�� ��n��M��f�F�AJ�Q�jhȢ���1?P(i!2��"Цx
�?��iAH���I�8���5�Y ��a�|�ƽ�O�:�5@;`2,�1.&�M�hh�_��ӿ>� ="	�I�#s��ʝ����������k[���ͮ����ɗ��Y��6(�_+Ps�zuW���k�y���H�'�v�����wN�z�7���5�5����ˬ˰I@�X��&˿G�(�4�0f%��O�#�e1���
G�3�w�8fU�Y�k�g�6��M��m4��'��L����*�G�F��|]��ߘ./�t8�:oYԾ_�`uRRleŋQec|2�=��W0����<&��"��t��I�؍�6>tk�����R�|�U���񧒣a֝�,�^���>_jo�͒��7�� ` :OiI����X�C��|�_>�$��$Ptl R/��л?=�;��g��*��5�
�UN�s(��w�*Ս��ΟU@����+��*G��)���Y�x��%vUލ�X�uS�"X�#'P�O��y�_�r6JB��7x�~b+�)⑰��&�G��[K���ק
f�<�'��N��y.R,�$bΧ��ʬ�o|�:�g`�v�
s�	 �wp��e���r6�Z<�	��34U�_/��2z:rl҉�F�ޗ0IAkv�̯a?�r�b�g@����i�	�j�N�N�?M���_��I�I�KD`Re����3�z���T�����H�@���
���i��G���������z"q���Hni��}�Z�G
�,��)[�=Vi*�W�Oc�*�j.����t.�V���,�t�a��
!7S������䕘�ƨ�5d��uX���y�]Tpd��LgA���`�:xgh Wm��n���g��kȹh������QX��+�I���a�kډg�z0���n-�Xډ��xOh���b��Sa�iz���s}�������l���8X�ZX�}u�<�mpT��监�w\p�Mi>��=R��I�R0��J"U�0,+ng��IT�FG���C��ɭi�i��%���r�9��\���
Ǧ�-<Ş���C}�~����f��|#@v%cBLS�� ��[P�����;� c��=���QS��_|ɓ"��A8��6H��X�^QH��t2�nn��װ��gp�V��Ν�<qh�J� O��FIH�T�<	6�`^-(X����v��V��>�����%�;K��Ò��t7w�DPn��[��ZF�[_�8�������H�\���ݘ��0�`ב x>�[�\�⸓�i���Q@#�C4���7Pk#x����F(	�/r��X�����ɽ���D�j�| ��k �z���c�$������yiܸzE",����h�C�����b�b���D*��.�������[]��\��]ӆӊ�{V�VN��0���5k�$��Ha~��s�ﬗ�ޘϐeW���r� 9}����f��i�vn�:T��in�R[kq��	�1i�|����ˤTN�O��U{u�!{A����w:���l�դ~LҒ��\�� }�!��|\�I��Y���$/�v���ԓ'O�񰱼��kK�Z7�H�W��$���G"�0B���]"Gg�ċ]�.X�;n��6R�{��Q�۬p����G�'��f��6�:�w-��@��>�)iii`m%�^$�\��Bx���I�ŉ�xE�������N����œ�h	�+�>�uJ��D�0�@�}�����]��}ݣ�k����%�A�5j�nq�oY�\��a��Z�8EE�q��u��E͚ C�TV���Y�S�҇'�I�,V$�2[�E:M�my�D&?7T�A#���;�� ����5E&���4����,�;�4�e��̦��
0��,2�v�|���ŕ(6,
��s0�E.�Ҡ�IX_'����9:1U1"[�ն5�;���_��R���u	�F;��uQA��������b��L�'�u�'^�����J�ƀ	se��?E럼!�>���r-�5E�]��h*���!��i�#4�ҟ%������YS����J$�=���'�L�Ȯ���SƏ�
��/.M>}��\��+nll��3�,�=<~�b}u�G�Z.}��0�}" �ɹU]vʹ&�����S�FK�<4���'�]�xXZ`�T��_4��sW�b�VE�2`�b�88{	�T�AS ��Q�����,�g�䔟ck�m��e���P�
m�.��|Gn�Cٰ���TTֈX_��"��'��"JӼ0�a�{25���6�Ȩ�_�2S�k�m4V�[[$c�� �[j�)�m��q���R�,�R��D.�.%{��b"��ݵc�M��_GiJv�j3`}Ȭ�s�T���ӮMz�wԏH�O���7�R�Jt���F"M4k^���b-��5�y�fk)?��Ł
y	��x�{:��V<�r��	�5�>�o�fH�T�H��^6i|{3�,�ɞ�CV����c�T�e�8a�c��d�>��Oi�.�9��=��d�Xt8ȫ	@��a����j��H����z�.`������!�Ҙ}��U�E�1�zfY$3��Ėё�Ƀq���#�'��@��I$��d�Lk�����`R<M	6�<R*�z�7��x���jM�iv�my�?���,�nJ{��Mk��|��0{�����4@�@M�8�������[/��Q_�~-�c�ӄ���OeB<�Y)�O��ǉ%��q�L$�)7�)�hm`��Hz�
�Z��#�/�g�zc�{=�B5k`Pky�ѡ i\߉8�t<��0 6|�G����s�X���E:�$8n//��Z�A��;�� $��Q�؊t�� �Y.�bk71��K��s$��#�s�A������W0����by���vS���.P�ό��~ rK�$RJ����C��e��\:�d��W-�r� $7��R��,��(.���re4�:.N�g��g� ΍��{����!޾�99��($f�Xl?j�Z�LR�t�m5�2��gk�ɗ?g��DJ�1 �Km�ȅ��j=.
�C�$�Q���z��m�C��b�a���D���T��)9�ڇ���Aޢȩ���� �b��B�s�髬G#>��ֽb-��1_�)fw��"�G���K7�< 5݊�-��6K/A���.�*�kTK2t�������K��W��Q^�@D;�L744d�dך���� {�B�$RH]�5���Q�cw�k1wP/��}̦l��Y7��� �!���.wAaasd��~�܉���5���Z�p19܄�������ȟ���Q�xc�����Ea�A!����-��3��r:2�}:B�O�p�qz� `\�Gр���TTk�Q|�N���E�e��j��}�#x���� =s�q�R2���	��!��w�:����#�y���Km��	;�/�a e�l��J�-�6[w̖�#�.�H�Bb̫^��gO��Y�PX�o����<�dl�������igC��` ���6�Y���"��{�7dz�K�GtN�ⰦR �w�R.�-<68s+fC��Bv����Q(@��_�re����}�kG{-^#μ�����9�Ug��y��I����B�����6���.@}��R�J����&��L��T�$�Te3o?����H�c�7�ˎ�v��թ���ї��кHd�FM(�� N:���_T΁���l_~�(�8�\KW"��H���D����l{:&S��pǾY�8���xq�}�P ��i�E1Щw���,��
��O�H�D��k1��V�`JN[�ً?�t�9T B�.�4=̃u�e~�G��u��	��'�Q�F�4�h�$�5��H�q���	��%�Z��g���u	V$�o�i�ȶ������ɔm`�D�����)��Пѕm���H���t2 �q����r�N��K�������=�BI�E�"�Ͳ�ȨPU�yՠ�i$RN��	@���j��h�yS9��~�b-�x��}���Z�J�ċ�ۦ��K��/N�3M/_��,�,X��',�dh�͏�}���[�@m���\�a�Sah�����{q���ĜQ���]��+�	 ��H��E����H+P��L|d$`��keJ��P�F�s�`ˇ�-��gP��t����\���R�>d:�9U ���Y����ר�N*�������A3���� _Aw+��0�FE�Ww1�r-���)է��2�E�M�/Lrn/�I� D�~���d�"+�ާ_���Қ�w��
A+��i�wI4Bd*��e�?^01���!�B?���P���X�B�� \����#�&��4qh�������,Yy��/qQ����k#o���[l��=�c������zY@��W��=b��~��b�`�L���'���v*\��C,X��-$�!!�/����?��K�wp� �R�kj"l����-ҹ7�f�A�(�%�#���6	_^��5��f�k��ɴ��s]�	�%�_�;��Ҍ�� �1��:s!�Ν;άe&Y�e��L����$����������9'b|���+�}�)	��ሺ8T��rnn��d�
<��)�e�h��|�	��G�}c?����]���Z�<��ZZ����\)5;��\��K�%$�4�����\���i�(`� �ce���0\)�I� ����?�gs�Y/��T?��j�F+EQn�۵�Ҏ�E��ac�g�Y#��b���Zkw�_/]��*
h���S� l�Dأ�<v��Nv`Kd�_W%��y���f�d?c�\]YI� #�^	����-K�av��K�B��p��-�_������-X�/Tm	� �)`�|66�&^@�����,T����G��2/���{�����ۥ3��W������Ȋ��[$�w�#s:���Z٨(�7�P"��w�~�n���A]�BY��sB��F��럺%{�h�P���p!��!��v�����8EY��nd[�.�
�z�4`���HDa���fw��e�L�* :�L5�f/���"2�� M��H�o@��D�,=�Ӫ���\���*y+u�p�v�N���CM�q%*���v�E~��M:�"A�b�����@� Ѹ����N�� Ye���"���^
������VL��� ��`K؎�a�K%kNo-���/�����Rs�~�o�v�����3-R�}����0��#��r�i���e�i$��k8����=;<����خ��W+V��>Cd�O�>���\i%ӵ��h��Adk�b>zע���"(��5��T�u��d�f�)~}F4C�#��)"���FsY+$Ҽ˩Э����Ъ�����e5��A�U��'�u�VCj�8��$���[99h U�J�A�,3��0���Z�M��m9�\K�L�]e ��]M7a�?��(J�c<`w�s��T+O�s�^XMi��g��?�S���-��~du��V�$�@�[�9 B�������^��%���H΄���<o��֒,+���~���J�L�U�ݻT,��+���؞��G*����Yv�]ߡ��ɲ�~�tځ���[s��5�j�	73�{�-i�(���P>�[�KMS_K?ӴWѥ�k��矠!��I�Ǳ�7J��8me:���pv
A!��]��2�	M--��C�nB�3K�>/Sai@��=מB��J��I$I�]����9�I�6qi�a��m\�_y]X*yrxC�?�T�$0ӄ��O%m���fAC����G�@Vo�a��gO6�e�Т7�8S)j�|��0��,>�~ z�c��r��k���ɰG�@UHA�b�=���OF�2��=��H7&�Z�"2�$�q�]� �G@0MJ7���]<~�7�teF��P��d.C�Lߘd������+��L����w%X��`�tg���}����L� �n��y��
�
�5���WVn�/����tӗ0O6S�O��9r���w�O���u����A~�2X�j�Gi��Z�(o��7_���D�����w��H��(�$���`��	�6U%�lR��[��T�;�k��-P盇!S��Hm��Y�W�1k�?�M��n�
ǁ}9�6�q)���+MM��2�;õ�y:
v��7� _q�k�'}V�c��,�kV:���]�]�P�_ld��ڽ�5�*6\�d�A�ö�(�"LL��9�F���-�Λ�(�f4�F`�e��^�Q:v/��trm�Y��`�	ɓ���d?���x��S���ט874	�5�]Q�i	��N�A-�R��*����t1a�7]Ry���yo��b�V����Q�1m���i��"B��A��ݾg�u�Ud��	�����pDc���!@�Hn^��_$��<��&��p"��)��(�����5VGZ�I�����A
}gT'����F��11��ͧk�m�N�׫F��4��I`
(&�0?X�Y��`-F�7���?3��n��(���< %�X�Qp�6���mM
܎�D�c�(lCo�}&���9c�ȍĆ�0�Ȩ�='%�eO�{����wf�z��y���î�j�F��&o��x�Z�zMP�6��'��[�w�t�(�BB@2��:�A0�v>;4)�8�H�I�8K�Ȉ�Ol�Ě���:��P�+��Z;$r�K�y��{����8l�6z���cn�~�{5+��`��'`���yo�	\��;\ó�"|��M���sd\�%d�;��~=�L{6eᰋ�x�4��,�����k�DH"�<iR�!�7Nb��;�x�5�s����a��Du��Y�Y&�1d���v����1ZE^��6�;���*��7�}�)v� �?�K1�yw��8gr������n��b_�֠���V��!�{1�ʊ��X��M~0�&˞� �S�;^��t
:O�{	�c�nƍå�y��/qLm< �� D��ôgh;m���V�����g����Z�"���v�ç�eN��D�n�8/�T�/��]K�/���x*� q�C��&:")����!�M�@y}?������G�ث{]�c���H�l�����ɵ������ɈL�)�t�C�+c���.5j��|z\)`���OC������c���+��C��?J�)ʌ�@���]�3�UΓ���o/�O���%���l�E�Ѷp)�,�ɜ��|�_W���'cX�YD�;eG~��Ću�0����0YѺK�s����Ǖ��MesU�QzD\�B��o����	}��1`�;���ՀCBҬw�����U(�ΐڣ�����?��Wǩ�Wkf�[<���C""��@���VN���h�����= ID`x��W�6�8c��{��Բ�;�7�=����LV��&y9��҉
D��YUl�����h~f�jg���~�sU�n�5� "{�a$67Ț�����uU ���7�E��;o'�̹����_}x������e�D�_2G��S���y�÷�[��>����`��n����rN��
w9C�}��9(vH�t�,��V�>NPX*Y� 	��W����XZ=t8�*\=���y�4�G�fu���e� ���5*�Z�Y�tl#\��5d�+Q��/����V��l�`ĸ�{�7lt]I��RU�f~�nտ<��0!Q��<��x�NF��� �ͱW����]�=��k5-������;����'��|L�(�m��p��j�^'������/���Z5Q Y�����=��1�/ꞃ�����{/���s�Ĭ���VDs-������{OZ� �T �vV���2��o�C���6.jj����%�t������XJ)�	�q����?�4����2�$iv�x���X�FxxlN|;M����������F2f�� \E�A���j�-�DI-�^�B��A�����	h*�Y�lx��A��	]�d7����g|�8Ju��rƩ{K"f[���TF���'	�HƓ Ti"�D �,�##���,|���ԛoO����و7-D��&�U���l`�'tt�y��\��A�*�$��]{5�� ���5h��	�"u����"?[��: !D���3�����@�Y)JhU2Su��� J"YHH�g�뷙^��Ei�U\u�F��B�>��ް��F��������j�1P�ғ�ّ�@/ʾ�g�b��>���bN<-
�����e;���S��Mi�,P��8�ͧ��n��ڮ��"Z�IxC�2.;���F��s�Sp�ǹ�i�k��'���y	�3��X�C���W�
���h��3��g��B���s��'슨Eٝ��g�W�T��ˉ"��~���L�,l		���#Z��uIS�Ep�O�������WeP��֤�����F�C�ܬՙ�]*�����e;�껡|G��w�%�S�w�Ş��pǏ��*�1�S�U;���(�����*HT�W5��+h��:�/u��D �M�[���T.A������pϭ�/n��{0(i+zx�>�[�������$��u3�}�q�XT�k4��M}�(�������4{GJ�X���a~o�n�ĎE�3�-�8Ne�j�*�_mg����>p���>(��L3|x-��f`����p!p��+'���N��x�{�M�$�=�~JC��^��4x�l'�/Ϧ^�eԎ���+(1��YQsγ�9�d 9v�*Ψ�A�n�P���8!�1���H����o�P{"�3����<э����޹�7-
a�^����\�;��DJ����E�B�G����;O
��w��FJ,,�~pdR�x�=O�����[� A�T�M�NlB�4e<�S���k�y0�#��+=3F ��)}���Ϛ�a)sNm_�lڑ`�Z�x�-`�/9� �[��l"׫���d��L�Լ��L�U�#�^��5��L��J9��
h'�iij�Ĺݣ$���q��tT���hJ�͡�n�.��ەq�5�Du���Qʭ����ak)�b�
5�y������*�5ۿ�����$Q�c0�P�M���^��.9�r^�����h7DLL,�����=�U�
E)?�i(!g�+p�UF:�oZ���Zp	����7�JˍRhk,T2��D	�mkk� ��oy���������E�c}���aC�d�&���aZ�q1%Эzgؗ���.+�ܩޙ2�{|�����}+Ľ�� Ǯz��q�;`��������zRB%���R�ͯ�r�=���9R�- �^a�o~�j��)͠E&F�/�f>�%�> N܅�_c4��B�"�cajg����-��ph�FʜR�_8�֋��+�:���ޝ�+��FY���qnY|�����=�V�)���;ĳ��+�����_�H/;�,	�￧4����ؿ���D�T�+n�=�W+���F
����=?�d�S<ـ�Fuv�"������Hq@�>g&��^o�Z&�/?���f�%'�Uٱ�e7TԚx?Kb;�+,�j'
����p=��eN�d<�w �S�E���$�Tn��6���J� {R.��Cvˢ�T��=��JXJ�J)u�u*����؛7@ϔ���LKB�J4�Ji?�.'���<`��-�S:j�Q��;NL�ƹ	W��s��WM)eyEC���3��W#y�t�cz�*x��6߃=��Cc�MD���5W�?���8[J�*�@K�˾���0C��Vh�x^��[�s�����p�	"��D�I���K�Q!�s��P6o�w[����3��)./�ͩI�~��cH[ʕ+V	R�>�xjݩ͊��
���dq������;����3t����d���v���8U�ک>�/���`����,�~�?�}������P�	 e$6lo�o	��io��K��H* e&d8R��f#�l�׺d5yn֙�߿��j����U'
���DW6,����SKU�m�'�4��U�`jF{�٬�#ǮJŶZ2KT�(A���r_��KB������o<������V�y$�-�FE@�.<�-��撐���r�Ox��aWZ��&��Gt��L���!U{��t�h����P p��ȡp���_S���#�<��X��e�ƩC�Cf���N8���ܕ3�y����o����a(<<�`5�1������j��>�A��j.�[U?�Ҫ���	��[�[���
��`4
���$�Vl�[4��j�v�ߊ����7m	�D�v�(K	�̻��l�-m��y��R��4)��)�Ӫ4��]�~FW��[7�1��N�8V/�=���Fr���EwP0L�R��R���t?����?�9�Հ��xR�D9�;6"��d̼Z�O�F�&t��q�|�ʵ����Q����`�y�d�ܨ<�+�=�պ����f����.��~ԭ�(4�������z0^�>C�Y�pB��� �����!έ�H�1�{/��h�2+�WX��*
'߃��P���_��}C�Ȉe	�爝 K�ɕ��j�H��!�����/w��l=�˸��&	X��
�f�>�>��-�Ů���حP������|�G[�� ��t�D����է�aw�} E/��)o�X�н���p�9$�%|��䩃BH&�s�#��D�=\�
�5�6=o����Ha��!H{�m���'T4�6� �.�DJ�qq����(w��N��Ib!�H}���W��[��� ���e �}���[S;�b!`���?{t�PbXFa��w�2䡅~-�52�v�l���������A]�ȳ���6l���� J��yL�90��5B0G˽v��DGGFbOaOb�+d������� D��ֽwd|��n�����`2���e��8�!�����T\N<��BZRxg�q��x>K�)_�z�P��ȼ��΋Ld��S���q�w���� ��~������U7f�Ǆ��X�{��Ndz�*|0���{�S�͕�%��+�`l�_���<ȆF͝��i���?c~?�pgaz׵4�(�ek����p(�jআ�.3��X��z&��Y1�W��^�|�'G�K��u��T�#
��.��7�8�p�hY�r��Ӟ�l��kY���}�19�o��K�F���OKK9$�I�H�ir�F�Q�Bt9����B/pl3;r���P�ذ�i:�sh��,u4Km�W5�f2���	a�ك��6MF���p,�d4�D����b�N �7$��\I��AK	͡s���%�z��@�6R�Y�'\� �ۡ�� ��Nף�F�,S�ᇺ��H%�t�n&6�������� E�~U��k?���lt0Uw��O�A�b؉p��Z��`���� ���|c����H�[/4�g<%-$��Z��۽��� ��J��0q�\�}2��s&Y�J�����9;M�{.�Dw��8)��$���+�peҭx�UXFȕV3�����f���䡝zc��|���RqP0H����X�~o'F��G|��]���nn��jľ,9!A�������o�}�i1�,dc?�B�="�7��\��H�~�#��d�A	���~�J˝�͉7Y�/��98W0�����c_y����~�{�Me�s)F�Nw|�=+��u͉��>��m��(^IN�=��U��D��F07%�V&Z?{,�ަ�"�{�}¡Ё�b��Oh2��p���j�C���m��RwښIz1�D�f��P�OB����ٜ/���s8����P^����l^ZZ����E)O]#x���`%�ñU&�+�o�uL�i�/�&5�VTS�8�D3#�L,�	Y��b@f����w�]��#I���sO�d!�����C���/��ۦ�V������~�l��gŇge�cā�{��tV<Y�V�S�w��w���LsPN#Efi���TN�]ܹL��v��f�kkKU}*mF�0��U��f�7&Ai���B%���yy#�K_��t�Nu����H��KWV�M�����	�ǭ?�$�6��_�et�A(!9���-"���ʟm;�vK��<1;胵c����!_:��
3R�q\a���d\*_�y�����M��s1�p�&��)�y�@�����`��� � }�V�ʒ��+�~,�A	�����/U9?A���n�_�)�v[���#��HB�^�Ë��_`�"��/�������2�8X��)���֑H��|O�:1�qLD��=��*��L�y����#I�&���X�=0o�J��/;R1s�Nns�fݰtc>z{� g�y�ʌ�3if�ʵi����61z�.����RM�rvN�?=��v0�:�
R�򝟨��T�LJЧ�-�a7�Z���LѨ�D4;�U14�bo�r��"���J�ce4Ɉy�P(~Q�a^�5�i�Ŕ�V<�0��ڸE�� �	�j����3�'�]�_���'��ڜYbh�ᬚ�L�lÏ���"�{)===6F�S�-p+49��>Z� �c�"�\���ߐ̜ۥ^���{��H
[þ��,�}�x��Wf\�n�X1�%�jr\�^ ��G�U
�MwG�Ś�e���Zd���t���Y��G�b�*�=��YqZ5qPkOf�v֮������:z#�{�(i�9at�E7Z%������e",�P����(i����V Q=G vo�
7�+1
�~y��U�Q|M#a�=�l�H�b�ᖞb�ɵN������b�^��Z���eO�wn���T]��#�1��%�@m�C��ʄ ��Ő�U`Im�yۣ�wj���=F��`��� W���\�.��/x8��%nt&ʪ�B�}�R���<*+�o�']I�PB�$���o������lH	����%9��.td"'b���I����ӏ�1�6-�{��9�t��`���wU����@\k�����a�ߘ����}�R��j�_�n5�߻m4=����	�
�w*hg���V��+��^��{\��\�G��lI	:�ؒI w�U�@lXf�3i�[LI�����\5�������a�}���M�/�9��R7V�QV	��$s?μۈ����!��lW���G�3�{�7����×��z�����X~��;��!3V�9�e�p����xL&��ʘ��t2&��ovt���L�Oi�2�c�*� 9����D�9ʈ&F����3U����4?pyT4
`*Ԏ>���]^i��a3�躂�������$�i�eؼ��5� 0�����sS�Y��,G����%Q��mLg�����ͽZߒHQ5�`���ȕ,K�����1F�&	V4`$2��k�}b>�c�+(E?'<�w���6�H�C&u �,P.�SheFDTT����  eS���Q�ۉKk�e�-�}���H(���v�8g��s��̲Y)�L1���~�Z?sR��*�����a (��uۓ�'}R�����OV ˞�]N��;o�/�U�7�V$ �"�I	b�1r�o��1Y�A��:0c��n�5*�hy�4���X�V1�⩵��)�iHd�Q�^�I�ߓ���̦p+���#�ޗ��Gs�#i�x�q�Y�N�r��Y�JP�vCj/��S�Kѵ� �v�8��:�x��t*팊Y�NL��mtT����wT�GN����X�o�J*'��B��R�o��_@t�Z�y�Z-��ksy�6+�G�����4ۗg(=P4W �+�W��/���BG��[viX�r	b�伿h�R?�o�T�'�rB6J�-
�@�$�:}1.��;n�)�L��sC��O���c��~��2�zKׁLw���W��ݶS�<�`���6'׊I$�b���Z����	�b�~�X��)-U^��/�xh��� �۔���"Z��=+|Yȹ���-4L^��*9Mm��6��{���W�� R٦��s�1Ȕ�P���y%F���#���R_�{���Wϼ��87#���G2��S�TDl������X|��E0Mt��}j4�n�����1��6��&�ؤ�<�g���D��矷�c�$�$�Y�Ԥ�+��Bt��)����;����cG0��_�'G")�A��%��"&��_�fv�+X}���ab�:[ؠx�D�&C%/g�dmvfr#�7�i���Ubl�*�Ք��Q�63h��O@i���sr� ?`� -��<d�٪:QvI�L1i����X�]���c�;��o��d	)�i����(O$�>n��({�����ғf�@��+G,��ʧb[o^���g/VD� �W��v�=RAW*Wp�C_��I���TU9�Ҫ���۫���;�}TK�m=�,�BSl��E�"1�"�R�	�iVBƭ�-�%��\�G:@2����q�nx�^�cG�b�\�&l��	��8��r�7;(M?�b�E�v������9�07��V1�J���uoPF�bo$Rj���J�k> �O2ި��0��ĝ����S�H��Y�Lt]���z�pmX `��D���$	�O�(	� ��m~�-jέ9��½�w))��?萇���_��h�{@�j�?�wTS[�.�9�=��5
*D@�[(
"(M��H'���(��
H	(H�^Gz�R�B	=���������q��~�x�=����lϜ{g��L�n�٘�@�/��"�O`m1O�f;Ύ���r�u������b��⽨�g����sV�]tH����_��s�
�8�wY�Q3���,�� 'n�� �'�9,Z�A-��I�
¤F-DےS�����1�}u�s��~���^Ǳ�[�����e�=�F�~y4g��[��۳@ً�>2x��Ϥ��Ҋ���7oR�,��]M�	}��Φ �|�FOR� g��U�ünۣ�����qZsk��h�Ѧ�i��X��-���%��W�1g߸��-�/p�����$����}J��8�G�.������gd�(<A���Z��As�d�X*��*`�1���[�.ݞ �B��#%nv�gά�uH�A�+3��P�k�����O'��&_���A��Km��k#�,0K@wR&�[@6�T�M5�`3�UϽ��D�/���J{HB�4�����Q��n
X K�t`^�k��5�@�t��z0&WU� ��*~�z��η��-{�H��vi%�T����A� Kp�t��8`I�:�f,L��%�3��#~z����aР�����7Dɞ��1��5�>��F�L��=�
h�4~{�·�۝�\e��]^$2��\� o��4	�k�Q �""Co\�2_F3���p97�z���*����C����/��*s��6�B� 1��lړm��5�l�0��(�>�Zl�'�韼��4��L����?���7���Z�1hQ��>����V�0(>�GK0�09������XuE)s� Pf�*�]Qq��d��B3�/:b555s@��1ϳn��8�r��3kޖ�b�20;��9N;��zވ����ϓ�+,%V����Ҋz�,�>��L���B u�dd�D�b��V���`���":�\u���M�� ���|e��b�/�]��$,�6j32tӠ����w�whvM7 ��Қ��R�K�� ���~���~��F
Itն������U���X���s�8v&b���A�H�#Yz���{Z�}�Wu�ں��U�����ҧ����)T�@2(w(,=�7��������n�	�����n� ���#p����Z�L򇒌�n�����f��E��@!&y����DZ�~�/�[ �$� �#ޒ\�;��f+'�35�K�K���`�gN�^�7��n�|B�UM o�ǩ�{E֮��a�c8�����\�`���ӹ��G�֓�������Ѝ�������7�
�V�Bu��7*4���p�hOТɫ �Y6��R����
�'�����I^dg��(C��n��~; �q��H04$D����m��
�22������i����p	��nRgg�+���휢���jv�j�k���z�Y���+����v��[�|�C!�
���Pɚ&S�i���nR׎�����Vf�2���9hw�I�m�#�=���Ô3㪐h]
�4����t. ���`�Qf$���#�`��H���Q�[r�T
9��f1�����/˰�V�r5��>��F/j�6�b1��KQ��E�'��,��95yݺ
:��n�&4�E�8��)u@W^>&�V�H�8�/��K��H�O��+ܕ@���)�[ W��k0n�kǗ�Sv~SWW�i	��uie��{=H�XX���:�_�Q�4��mCG��K�3����L24PK�Ȑ��F���kY�"Bc% ?h��.?��$� !''x*�E�x�q��e!p��&X��7���(�1���R�H��h��eZb��&�u�k���������7��US�K^ML���p5�\ݒ�U�>����S9��A�����3���a�~cZR�Ǐ *w��r����[k�m7F�pC���@����^t�W�hT?{a0�Ǧ�K�KTO[u�qp��m"�: |}@R��Ww&��.&�Fy�P2�)h�͍�"\,������#���PE��
���9��[�<�[�3�x8���3�$����j�Z�-|��w�a�k&˷��jU��hU���{h�<��	-�����$E�!�E���9������n�W���cj�"���$�o���`�c���+�'�*�,q�n���ļ�b��ǧ;d��[�)�+��Y��$G��e�r�����}T� Ց�%�ٱ�.�Pӎ�ã<�f�Vn'�Ww���W�f6]��R�4G�[6~҇�s��vôS�p�
���k�O�V�*~�I�����d�����&�#�.	�6ם*�j� ����Ama�H�eR:�R׋����<��F��
�:�?O����P�AË�T���+5c���-J`��+BI�dS�����Z��<^\8Y��٣��TMM��Tm�	�	;�d��Ŝ£��f�b���@�KPQ����$#u�\mӓ�S�<5#*T�U3��S����%	~>R�)�v����"�����e�x�
i����X��H��v�:i~�@��95j���?�f'����V��S�?̩�7�U���RA��&��El��P�{Y?َ�/?��ѭ�v��j?αRe"�2Q�f?e��(��~�A�U*��l���]��Z�VX������� �����RO�z|h���l����O����Y��N�IkG}ۓ��d�t@B�4g��tm*\�u=��O=������*�����z|CP�e����A�R����T�� ����.�kƹV�hΰ�l�,oY������Й9"��W=*@�z���9X�s*���X�)�-df�����'�/8��T]T��|��|�C�!BǏ���h�����<Ԡ>��u�\l���yúQfX�T�VT�\_� �T!C�8�c�n���>":���S1ڭA��g�����h�.#�1�H�n`�1,�g}��E{��DL������9q� ��
�s0�Q�����tY�\`T�a������OoS�Z�+zJr6xxG']���t��g�l{����UH�+L�Z������I�*.�j�V~���
��R{:��~~���#~�0�,/U
�w��-1��Q����^F���⦵�c�Z��û���=�{�6�� I/&M�;r�1���
�9�FU�&a�<;rgbD�`�1
I��}	d5è���I	��$���}� �����[�f"�|���O݈�n>��DvP��((#�1)��G�����.:�'���-X��,�h�b?�$>����:B���h����8���VE�ߡ2�����Px�45�W#�<��¢�e�6�p�PO&�8� ���;�^`��l{�jFur�P+!@����c�d�=�P����Z�3,}��h�:ի�in���Ɲъ�	��?9�JL���wjO��iL1����O8?��vrN:�9T>4�A�v`�{�^�
��%G�^�ގdo}�\��~c$�]�:���k�j:��tY?��-�zδE���i���s�j��UN�$R�U�A�h�^�0��K���[yB�.K�g0R�lfZb����}�۫7Y����+������L^�d�U�)�E>�\�ں�1r�vB�*��HeJR9�
��/� ���P�.�J[�Ti��j����0	����UV>��m?P�|�����5e���������j�(	+;B��� �S�=i�::_
��H%Q�5,6a�	�Q���ѝ���%ahȥ{;ԩ��An�c�����E	����Y�s�Y�%�Ws%�yb��ˏP�㫏W�OX��/ϗZ�焮�-��.52�ϻ�i�'��w{��-���qH]=�k���Po�G�k�l��'�Sb��\����%�& I��"���,��^�nJSY���'��c��DdA�(�,"ɐ��"��^��C7h��zW45}֍9M��Л����IG���'l��d�u�����4��]C�R�Ϣ����� ���A��$���t"�-S;����,g�SJ)�::}�4���S���m�����B6W�4��K�ȷVb���]�T��9� z1!iE�Mܼ�'��1hj�3I��j��?7�.�F���U*%>�X2 |d+	�g^��]O��O��n���s�ǓHǝی��Ʈ�R�uh�g�I	��3.?I���B�V?'���'����&&s��+d;��kx�9��w����e.�='߂�hC���+����ь�M|���)d
h�2�����/u6_詹4xI-�	k�m�s�]�_���֙T��]��g;�xs ��ޣ�����)��$ �̈XC�3V���.K}Olt{'c����\Nu}�%+�n0#f�?��T϶�̮&�6�s����N�n��,c'�/?���j�D�Y�	�ʯS�����Sོ��"W;��C]a��r)���3T�v��Lk#ߓaO�.�4��tk�u5���(Kܲ]��Qû�e,��Q�q	��N���v��nn����d9�D��\X"�v��Gt�~����X+0�>��mѴ}���Qƃ�.�]��8��'����ﱖy~��.�԰m��ڇb��P��W�9Ƭw�^[5u����SexhZ���Y�Rpj���W��Y|�%�\��(���i���.�����O;�c�s4'��߭ �W3����E(k��a#A�	�D��c޻�K�|A��Z���l�U5:�м�����F���]�f��sgk]m�Cx�H�A�M�������\�b�Y7��D/��k�����~%���z�|M���&��ߩ�Pɪ�����mC49VH�2�$P�HX� ?��=cɯ�q;��koT�<�$u���*�8����J=�؍��,p����)M4�5�~��9�h��C�"9;.,�J�:�[n,	Ȫ�%F"DO�?QcrGN������n(�'�{͓h?}%⁪[F2��y�����$a��sI$~�V[�����������[I�y��E��/M& ШR @hUBB���V�U��_�,ñ��Y}[|`#u��lI!�xϤꣾD����ѵ�1N��B߁�`7�*0b�?)��Q�?���V*Ur��o;������&��6�nx�W������~%���q�r�g����}`$�L}��^|������s��E��}�T5؞��䒗��i٣1bAەx}�E�;����c�B��I!��jHMBI	�q�$�p�݉=>�.G��O
|���9�0���wB�� |��IVRn��1q��O���(��GzSS�ߑ��\Y	'��1e��G��T�Y<3�,�E±g�����S�U�.�����VQ��?�>3=����2�O�I�\��27z/�����퇰��	�I����@tl�}�f�<Y(�$��H���C}���М'bߋ�w���p�l��H|=i!��B�O��JlFT��
���!}a��w^v,�
�����adݷJa���uy��_��yw��3��H���׮�Ɨ�,tܥ���������8��ɲ?]�SD�b��O����'����_���O�	���>���K21雔��[�G L})�_�h�C�K7-#FQ�Bydl����ձI��p���X9r�^A!i�>�&l�󱦻ڇ���[�Kuaj ������\Q�Ln�˱�uhU]��RՀ~ f���c�CjK-L$�б��L������Mu����r�y��8O�� ���0���ϭEWpy�Q�V�p�bg�o��/B��,�<��U���z���L>���P%��/<�`a(���ᾅ��L�p�*Oĸ� �ơkR����O���&Y�W���䩀P��ꌹvP�q]�BR���AgJ7����#�4�'����-	;�0ə��)z��9��f���	9��Y3�k�KmZ���jRީZ��.7���gXQ�a����u1R}}b�"�KY�U)>�_�X�u�b�����KI���d��M��uRO�Їf[khXu� ����">�%6�Ay�$���p��`�t4^������+���]kd�n�x�%6���&�?�����UT R<l�jEz��^���x߷��by�j���O$��|���ގ�	���26e��9���rΑA�_RGC�4��۽/h�U�~��E4N��$�À~�/`\���� �W�ǽ��TE~yPƯ�2��]@������W���
�����(��W]���(�����rH�����ĐT��f�����R�=|.Y��e�,�4��O���8�8)t�Ƈ����+Z[4����ꨁ?>�D$>� Ѡ^��Rkvw�q�i;_
������W^��ii	g���O,V�=��R���Nrs?y355�'��א�]^���%��%4i7W��KUX�g�dgn2ִ��x93W�
K��(��LDڟ�<�V��2�Q�
�A4j�-a�����ȗ*F]�0匈�AnJ}Ή�֔h�[���b�9io rF$�U���yRO����Zݛ	����p���mHn�,�~ms_Q�?���5��ncoxwC����4�Js^�>S���E�l��#�d1L���Uk.U䬭�Ʋ�V�Q������D�����ƿ s�	Y�hzY����
�C��;�I�0Ǔ�g��
�ދ�������_lJoj����+��5{zd���}���w�P�u��/���	�X6r��2���wW&��"z��CS��matt�� _zx<%R"L۴�nҟ/��`�K����~]��y�V�H�v��䮏�q���@����=>vQ1�J�b��"$�6���#9�N�*���9)�IP�1O���	0�wrs��/k�cs��;�]��,V�;;Re�Ml| }(o�oh�2� C��k1�c�`���K��wk5�[��^�4>j�][6��8��t:G�io�f�'�C�Ѽm��t�������3�c͡�𕀋����6ѱ:��W9n`k�p��7�HA�6*ʾw���J��4^�[@re1�������)/�U�~6��s�d�^C.X?�S� 'Yu6�{��=���^ޕ ��u�Nz��b�Pᇔ����^�{��9�����Ǿ���������kJX_$�P�����0�^[�f�pQP9�3*ok���0��FZ�N[����]�C��z����9A:�*��t��>�B!ij���x����<�N��ǎ��l>o�1��\t�����6
��?�����
?Œ:�o���[W^����װ��+'��F�%N^�Zu��k���:����P�6�P��=���K9���
^gx�[V\ҟW��^x�Ԛ�%j�;'���C���q��.����1K�*��o�'8����Ú�>�5)>��$�;��ܧ;3<+����V�2�سp.6�I���w��r;*��DL�(����]��2yz�@:�7ɍ"!���u��U7'�t]fbr�=K���!r[䑳˃��w�>�fhA���j+S�Ǒ�
Φ'[����<�Q�(�<Zc/A� ��8=��Jo�y��J�od�W��%z]ɽ8��3*�w�g͝�F;�2�d����-���t̧]�	:4�QΡ���;��R�&�
e�`��4g(�W�{�&�n�(���F+$&[�m�S�|YA*M�=f���U�D{$wN�*Q��O�Jw�+��o�N��6t	��s�N*M]�o��㩶���#���q��▬z�א�ɻ���Ճɘ>Ҳju�.a�v��me,�=��CD�\���kd�8F,�"�LQ���B4}��6�$���qV.yw��p$���T*�S���䗍mA\�{�`��gP�v��P�L��*q1cl�P����yF��-ʊZ+�sn�+����(5���<Q7��_�H+��C�2*>k�R�Vn�%�r�5U�L��W��ԦV=I_��y��|B*���l���"��Ҡ�B���
��J�>狹i���O��TGcG�v�a�on%j����z1fk���@+���Ɖe�@����������>�&����D�^k��x�3�SIPH�n���NU%��BjОd�p��\`�2�`UP.�u���jP{�]S�N!ӂ�\".N!��Y n��V����=���D$Y�>B�}�>�J3��'��/T�]�KP� M�-0��J�$��<?�K����j!��E���ڞ��^ǭ޻������A�5q����i}���^ͬ�F�|c�f�ω'��Z��w"�Y���:3��h�4m�H.)�R39Y��u�T*Te��ګ�P���T5����<�X �̃Z��$JИ�E#�㳫�����	/�x��-W
�KCJ������{�e�a�����n���y�d���<p���z����f�� �:́0������ �}�D��`���F�PԮ��L>��0D8a�\�y<g��e�h�f��?��T�%|�8�2���5�y�_�VtiB�v�r?6ʀÔ�ѿ��d\��jy���ڟ���ȭ�P6�F+�١>��.�ݥ��;V��%��������
��AC[��I�@[����¶Y�ĳ���t���:�����&]��H�T$��9+(�|muD��Df]�V�]�K����P��>d��0�[֗=�|��ZXi�P:�܊0@8�CM5�=�휎<n�A�x"�:=PT����1��ܪ��	/DfI!
UY;�K��yy��5��W�m��1�3ߑ9N���?�(">��LɫUiA���Q]p*�(T׫�S+ז'������(?���w��K� U�h~�e�.N�6�C�9��K�P���T���p�V��k���vC�|�xC-���;��׳th��K���$^�y8-U�YW��L+o�l;��.�ڪ��J ���o4N%�����7@,����q��~��H��G�s���8Q{����ar��ҭ�ϓ
{Ctdܯ�D&{
���#��/k]p����	;�r�7�@' L_T�Os*#	��K����:���4���.��=�Ჲ���J��k����Wx�e3_8���W�;Aז���m7��@�/�%} ��qA
"��	d��_��d ��m�kc��/�yyｯݬ���f{�#4��´����|_��b�Ԅ���썄6q�&��O�T_*<�{:��I�]��]�yk�
o���Q��8�=t璠��S�ow��w��w�n��~\���!��O]�#*��hq-���8�D�C�G�q|�Og6����v�����@�{�;R�x�lŃ�/L�v"d��S�.<�y���g6f�^1���;�E~A�~�%�s!�#U6^��'�˲����U:)M�u��La�fY���k,vU���:n�5�U�����H!����M6�{A�.j���ƫh�g~F��&�k�	؁����)���˽/���b������o�Y�̚����˫hm��������.9دeIn.�F��oьY�r�Q���T���K�3�2�x�-�oJ�O��)�)h(#MCK�+6j�y��O��h�0�뭱T�w~�%�Ծl_�j��8���'���a��U40�!��ܢ��5�����j��EQn^m��Ŏ�bi��`K��CCǥ[��l���)9oCt��L�L�!�v�4kxa�4ܻ����X1�(�YU<����O�
�^�s�C(JkGjX8��d� �[�)�5jiU����ߓ;�_�7�۰1	��(M�76�4mё_$u\Χ�Q�#�&��"�#��_�LY�_	x�������\+�OϿ,����G=�l�բ���@{��+��c�O t�b���涮S� [��K�L�e��|f��{b�q��$�eڀ,���p��n`���`�
�]�
`t�fփfE��!ǋ���7��ц���:t$��~�;�F��-CMSծ��X������ǊuT�_�c^��I�FXu��b}!ڽI����Yk�VFUD�Fl@��Mٰ���k����)�S��6�����>��ᯜe��i�b*�CV�/]��+Jpu�%م.�ڦ��K�Ӊa�7�M1 �L��g &
0��9�-+��S+��Q�&J��㗍����ߧ%�~m��*@�/D�a�z���"�y\�X2�Ok�fQ��7�jB4�[�s�ۚ2��k�r,��t�usJ>�34b^VuLu-�*y�c��W<tyʪ0d8�`�٫��Ĝ�2�;��{z!n��P���c��Ȩ�o}�]{䊚�h $s|`M�R��i+M�����3}���o�%���=�v�M�iŕ\�SV�>?ZL�oY`D-����k9n뙈zG�k�V4���K>ܫ:`�]����5_��=hC��s�Z�Ɣ�y��ŔX�e�Fs�	pV��0�w=�ۥ�@��Y�SE��a�I�&�i!ǜ����n]KXy>\s�ch2�Ϯ�ޡk�1WL.��5�λ����<@�uE�0�Xpۉ����Fv(,P-�@��".\�����\��ܼ��%�<�X1�W*>�C���f�'�n�߽����<P�{ ��[]&
ľ4���A�[y�XP�Lz��XJ�����fu��2�M(ׅ5�A�8J=��n��{-55����[[�����z�J��Jj5�D��+���P�dQ������h�5����"�a-	6+�"�UHTm���Y�y��u�FS����v��<�b9��=v�ѡ=љv&b�q^�I&MZ�0_ւи���XT��e{��5��aA��>� )͸����V��v��go�jD,�� pH1Z�L3�Y׼l�<@Jս.��`z�*�hJ�I�������|��E�I����`�$���w��ڡ��\<��6���}�غ���sA�'$���!=���2o�|	���95��һ!ȕёb�}��Ux!�f�e#J�}`
�O��+��"�z�N���N�θ^cb�)�|�E����Um٨�[B�"���-��))_����f_�3�漄��w�n�c�,�3�vN�x�(�-Ξ�9�"0��e����F���;7��?F�L1� �6����X�YhO K�Z3!�..LK9���g��A���[Q���|��\�#��,w�H����ۿ��ލ����m�1�}y�mÛ$&��q�q�:��8	Hҹ�j���F#T��⥜r���ue_i���8v+�vt��S��8=�U}#Pu�u0^Г��_-�=��*밼�����N�f���Р].\Oy.h ��s�P�h��W�����Eg7O!�}�>
sk��pZ��#ﵬvg�o�����htg�[�G[�|M8j�9��gby��A��������Қ�Fc8t��3/��U�(��/�X�U�5+�R�ǃ6�>�����N��ɫ�斖� �&ే&��4��@�[4���X�-r��+������Bl4c����	�X(�r|kmߴ��pZ�ޣ�zg:h7��\gem���&GGϜ��v��?9HH�n1]�dV�*�o� � @@���+�Wt9�^L[U�KB3�u�Gvyh��-4Ꮚd�T������Լ;[W�fX�(�ƣ���F�k�z5B�TFUFO"j��#�e���-��`����Y�o|]ׇ@��{����ަ�Ym��
cNIM� p�q{�ln����v�85el�RP��$ �<���u�!d�$���HO��44��o���U��+^����Z֟��;;��ywi&[��m�Kx��G��8��ӗ���R�X�9Yd8�����g竑OX%�D�Fɉ�+�.�T%pY�i�;�4�CT�U4�$|������v琔���J'���ͭ�7?�fЭ#U�x/��-Z�X�Xi$�����v��֭�Ĳ�'�"2J2,Hs��hT��|҅FJNMM�:a}��Q���� �[\\�1Z^�d���ǘ`1�! �o����'���y�I�k��j�f(�Ccs����ZG�J{�YE"i�����%B�9Y��0O�]��J�>mh���y�����`O��4��Y#��xs癱���v�C���9Rr��v:s�Wʶz�z8�N�DI��y���snD��+x!kr��&�Jkh>1���tΜ��7ă��E����өa$>���m8��f!n�����t�Rn;��@���iGb�9K�ݡ�Ϳ�%��l5l�mN
�+/^�F��rZ������4�#��}E'� ��\��&S'��n�y��lN��Z=?�����cY��X��� �IAN=	EW)�G %�BkP����P0�ۤ�u������'@�+�v�lg��*c��F{h�p�{��u/_r�a<ދ)'�X@�I�����U�����]�n�2򜎔�+{W({�N,�Dj����O���B�����H�qJ�4耓�:<@S���f����/^\���Hx �e��ܱ�'-��Íh��H�M����[Z�F�2�۾`�]f.8��m&�ݭO�i�̖>���ѓ��ޝ5�͚ͅ��ꐎ�]��A�ɓ��-�8�=;;�?������*(�/9`@�<]�Y>bٻ����=Z��� 	S�TU���!�:Kĩ�����9`�ڻ���@�oO�VK��v� ٹT�r��g���0��|�j�~v� ��a;��\���.y�,���6��?�`��:__	u�5c�D�G�}���Yt��T�$VC�r�'�F�l螬�[�nS�B)� :�!#%�+��e����� 1�.~��=-�6)z�Mk� 'X�Te=;@�a����	���˫k�x􆕫�{�n�~9����G}��<�6$,�f�	WZ[%��׹��\�^c�z�|�)��S�����x�Hm�����[$]z���Bl��p�R9��x_�sV�Ӥ��i|�]�щ�OZm�[����U�Zz�Ǐ�)�������n�*j�� ����m�R�����66�ݼ���S���Y�s1׳o�QF�s݇6����y{+����)D���s�/+P� �N������K��:^O�A}P���ꀏ�ޯ����޼�]���F��etg����GG�u_u�Qd^YY�zIC���g��� g����.l]�Fo����#����hWӸ��ǝ�;�$��?�S�\O�yVn8Ja2>PefͰ�\e)9�(˸��8�D���j�azz�
�E�-4�Jtn��Q��]��G�"g��$�?�@�s̺���?����/�xu���:8��S���|(ݥ"_�m�qR���	͸���
M��:,�v��3�QA�|���P�4�\4A�h�{�w�;�;j�]�47��.��X�e5�40NْS��U*����΄꥗q//a�XB�lx�X>�O%���|g�@��Y�\��=�{"fD��G�΀bM+�%���W�dS�ʕ�8z-��9Փm
��.mkm�~<��0�1]z�Fd��_��~s�*�#���B'����~��\::���I(W�+X@R
�jWjOAA_�RE�'5�w�*q����Țz���]�%����1M����7��[��s�[>����k�{:2ǄsH;J���"JmO�(W�'O����TSR�HsDڕ6'Q�Hך�Y�5�l.j��$����<:򮾈Nm_������O��T����0�0B:�$��[�E0���r�$�mz�pIIiR&����M���iڙ�~��W?����/ƆC���S����H��%-�)%+�
��K��U�is��ϊZ�X��q۹��&ݬCCC��w��ĳ��?wa��W�{��Z'�1����y��THGW#]��vM$�����6�Ji����
e���T��a(X���E�(�n:0��{P�����+"��g�6���@W�IU8ûg�1ѷ9:e�cf΢+�K�'�6�%"]��띢Lq������Z�H�EHx�؂�u��՛$;}թ���\A�S[>Y�[X��6����' K�t����W����Pz�P�.��T@��������+�,�R����ޑ�\�=׉=3Y�M�w%V�~�gs��Sj��O�Н��W�������X
z}�DA�V��"Q��g9�� �OǦ��s�ͣ��#>�֒���í�'b����{�}/����E�`bo>:|B���ρ�/�k�կ-.oV���SQ�ÿK�K���P�n)�It�P���ĺo<}�)IW�V;$h5m�����z)3��>�۩���C��8��s+XI�5cB�W�*U��/l������ze����k[��Eih�;n�vj���ߕ;Gm�$���-���u>���������s�~��y����p����� �8T"��!���7��?[���}��/�`��g;�9��-���Ō�|��k[;}C���O6�,\��iYJc���x-��j��������龧��U���
u��z.�8���'��p����%˜��`�{��K��-Z�y��ȇ�UznMY^G�&�yl���E�R��X�4���w�·��Α�`�A��8��fjE
t�.�}n��xFz4�������L�NE+��$�W��IC������\�j4>	�e��y�ݬԽ|�`-��1�s�d<������v1A��k��~����xJc�uYɃ�Ur"���%.8��@���90�g�D6]�*"8*Qhl#�����Xln���m�Xf�֩n�k��&���{N���ͫ3+��k&f��>B�&&E+�Sʓ�$�0�$&��(���ǯ����L
SfR�*���H��ERP3+���K�0ԇ^C�� �1'��K�#�MMM�3s���D�&=�i����?�^ЗyB���	�-*2��^]u��}���_��6c)�x���
_oŊ�T����&��X�����Sv�;|�?��W?��ϙ���_���_\��W׽�	IY�MbFb�����{�hZ��Ueܶe=��:G�C�z�d	[�Vcs�,Y;��l9?$
*�?��o�ϗ�����S�[�u�`+׹�\P�ӑ�N���b6�er_a;��#�ݺ�r��5����~��G�D��UV��6�~}��b�
n^e_%멃��4�^��z����Q���E�9� ˮ׆�Q�Ha�Q�K���:g�d���du�/e�׃\�/���[�M�C�V����;����ʾ�eԚmj��%�?Q)J��h�#��O����EM/�(%�J<��[e�ᢰ�֞�׾�*Ŕ�����d��-��?�P�f�i�6j���?�L��ea�fev{}�=������n�3R���y�[���n��kf{O���}3��;3">*D=ݶha<���_��>��9�
�l+((HZ�g�Z��j��>�m�%h�p�6Q��c}y�l׺�5AF�o,�B���#_�yv~�~H���?����vw�:F}�J�@��I��9�^���〇���$����r�٥�s�Qc�%��I����!;'~W0��UDe���ͽĆ��ӓ�QV��
�d#<�'�y3MJ�^�R���t��������}9J94�~�t��#��.��C$�3������g��nf��R�R�G��u�r��9f�F(Ok~.?�!�[oůlp~�������x|C�����Y��.�����=�uO�	������P������'�&�⻬m̈�sQJ�t���ݹ�I;}v?���?��?"�#���H�)zg���ݾpH��jS�1K ��V�P��=Hw�l6�O]1J��He��Z=2���tj���{κ�ǟ��7�v+ܔ-�BW[?��+'I���X��'�׼��>��9f��:�m�Aw|�x2�d.�`V��ĥA�យ�(�@_�%���.��,"�'�o�s�I�;0�[���1�y>�6oQ�U%���.���[�C�t�C�=�[dm��E)��-��#�*{�֖|(�L救�xUS����$�_�P8���[�;���iѩ˧'�Ӷ*ػPiB���'�-�|;�C���-�2��t�`prk��1��@�I�>�C�a~����k}�)om����v����Ob�P��דs�`\MIXw9w��6���#�K����&==�[s@w�,�U�9n0$�V\Μs�ۓ�{�b@1�[��?R�c����*u�OJ꘿��6+�El��۬�=@*W���҈����O����DY��y�Ċ��ʷ�����x�Ͱ{s����F*b�n]�����PtVn�+�9�����Ğ��S��rW���}~E�_�$+Vl{X�\w㪼�����xM��0"Xtu�b'�����z�uM��z��#V�>B��&�:)���ZZ��/<����D,�Dqf�ZJƅ���)��6C*�x�gVz�����Yԛ[������}�oH���=�A�G[/��8u�/�ۓ��ƶ�+������ ��]�|g�*y/�_K'`:�WfV����׉�a��P㇎����e�o����Q�S�R��(�

{����t��-iZny<R|�����Eov&�I�������.M<��6�n"
(i��?���9�����"G�}�[=e�8�Bt1ia�ma8�ͅ��\�F�_�v�z���ˇ�_:n#�O��S��s���Bh�[R��?m��:��o�?NH9!��Meke�ez�2�+6ce&��bg�3⳽��+�Ҍ��R�k�$/���~97��J�����߸�Е�s��L�������MGRz���~���vP�v����������)2A$�ӑ�n�ª����N5����r�����o{׸2�AŻ�I���tmy�O{�<�m-nxm*�#�,%�VUs�u1�_����>��U�V,:��=��ȱ��q,���_2<�"�V��#���#m.d3�:��Y^馻,tt�S�itt��=JV)�r�u��(=5�r>���C#L-����&߭�?�m��KܹKmh'�6,�sN�H����ҝ�m����{\T�Ua���������Gz)��u�D�
�?zq��Um#���N�kV>�g�Pm{%������%ir���b���f���C�|��J���׹�+U�m�v�6�Y�K���N�n%R�+�K��JS���Q����R�Dr,8�'ń�0��e��D�bj�*+	�&��2�������&x/�jdk����ֻU1��7ݼf6�[!�m���z]����C�����_#?��F���Iz�P�ܩ�j��C8vc���-o�EX�EU2}\6cd#"�w�%|�N�ן�������w�W��bB���޽?�;� �N�h��UYZ��������EM� ���թ�����_���AOؔQ���gO�~�wArT���MV,ݫ�W���,��(����<v�O�ɑ/K�w��)����I��E�t'��d4�"u��Q�1(�[hq��/6�ƴ��|���cbC�犍��8{_M�eդnz�L�A�a��� oL�K�.���Zn!��d3�_�(�0������_p�i0��;iӚ�!R�l�6j�༉�uH����ߗ�.���e9���u�%Ň[rž|S���%��~1Օ��{s���kf��sk��P�0aD���2_���/O�}�cYW7�z���J�(���e��K�ߑW���c7>n8��>��;}�|�G�]���;��.�[��O�������?��
�E'I�$9v)G�.��f�k�<u� �[Ju���q������Ys�VT�[H�Sf�to��i�P��/�9'Y��K��Ysi2�r���ٔ�]=rcX�.�9�)�\�L3BL��?��;���}���bAQ�bDE�"$4E�w�
� %��F���HPZ��!�"EP�z�PB�3W ��;��s�8����1₵�|��>�\s��|{f1��xx�3�|��x���3|O�iG�B�8�m���r�'�H�PG�ʱ۞�.I��Q��W�?�[+�&�Rb�`��+%�rK�x��}�_��.)ﯖ�A�9tj�̂肏�F㵂��y����1�4���O�,�J/.b�H�btuS\�\r�aolұ�q�艜�������`0U�T]R����R��N`�!���	�g�	i��jfƹHV_�6:�]~��z�3�2�g��GI nqR�#�Qg�2��C�2c�b���u
�eA
'��U4���eϸ-'|����E��+������?��/�k�?�D*c��[����ѥ���c�u=�Y���R���C�t� ��4���7$Q��J]Ӏ�6��)&a?]�d��`e�%/��.g�5fae�Dc,G+��~!A�2	-I�����r��������hJCʺYp����C��o�S��U�I�A�J C�E�^��/¨p�˅�.��u`��**P ?"z�/-2s!�y_���qE���ɶ��aݜoB��:bhQO֍�ṷ�A)�S��"����,�E4��;5�;Yr{�������dN$r��<� �%���K�i���N6d��w�}��x;�޹v�J)�Oo��q���h���~e4�P3��� 1�;PhL���F�j7�$Иk�loT�h(&�Ԥ���}O�g�ꨪ+��} ؑ���I��Q&��Oe犥���bG�mV���w4R���]꩞H��p,~;���q9����O]3^����R6���i@��<r�y��,�RW�
����:������G�{�vkn@�}8���*d�G��%t�[M4���0���xO{��<�IYf���#RE��u)�O�2��Q��o4�尿�%6�#�֭���>HJ�����
I/m����s�ט�s�1ӑ�|"D�U�˺
��(n�TF�7]��`���N�z�7i(���Sq�ֵs���X��҃���׿���{�K��K//,g�:j�1y` h��/��r4K�r�PM���m4~Fc�GISQF�㸨kB:�}�;�/@)ʛ��&fd��0����e�
�**ǷL��{+���x��8�h,,sA�=Sc;i�����#�&����J�W����#��U��0���n�y��V���N��w`x��6&��p#�i��z��<����*oi�o���_�w�_4A=������>"�^{��/vG���/���b_!����M`����+a�]��_Oz_��y��"�]�Sxy��G�������'"�Ul~3:!��+0rCc��R�N�7�r�/�T�r�&���T�괛�~��0����C�J�h�oZ�l��w�,��/���2χ�p�ع]��E��^��jcS��jR[ӄ�9�lK 6��.GT�l����v�1�N���R�g��չ̸��	 �_t�U�����,�7��Td�{�zg�#y�0���S��7�_���o�8�
���� �h�W����<弴�Y�R4kP�h����@f	D��=IIzq�ɋ#�_�P����6��2��
���W]����_��7�t�C�7�u��+�h����;�N�dN��?����@���F䩈Aޱ/���������|�f�ς��l��3B��~�ȋ!(�v�<[�D�n���AvW�/{��V�W����@C�<��y:C�3Q�2
�Q�"�So���=Gt�ܗ��2B���Z.��� T}����B����&�<��V��";��?c�4� �bW�]Ruv��Ի)��������ޓZ���IR�h"��g��^��?P���Q�ʗ�O����o�� 1���"R�_d����q�S�i�uɢ�{������N~�}�"�Z�X��W��u�Cc����{��-C��9�2ۍ�OǈK�e��}��\ 
�l�'/*ۊ�ك��w���&(G��[H�u�t���Ŧy�{�L�by��,���b��x�\�jSE*u�Rn��
��xI1������}"쾖@�U"r����A�=R0D�X��M/�$R���ݳ+ٓ 8�d[��d[j�}����#��T��^`ey�1(&!����9��2�H>Ewz��X�-M�tK����Oɇ����d��LN_p�Zv���v�nn!��ñ���^	��J �@a��Δj/�Z�V��j��8�~.]?���:�V$���)�Y3�l�a@Nk��$�r�z�a |Dws��zv��r�cs�g�
��oQ��J!3���K��+g���Q�]���oZ�[{�� ����{���M�s��|��\'~�݄v��'�Jy(����Uc��e���i����_db��B!�;sW�{�v���x����5�aU��2�}�&������Pz˩��� ����۾*oh�]{p�co��z?
�;��IC=�	��	������ {����Z7
�Fr��뤘'Lh	����fC .c�DQB�Tcm�'����'N[�LD%&���
SĔo{��k��>�9=�0u��JWJ�eI��=��z}@����Hr��Ձ
5��8��c����4�c�/,J5�A	wk�����Gd��9���� 
�Ի/�%�@q����2t��=�󏦅����f�8��Hl�&��n��.OWX���s]UV��^���9�z�z��~�F%����IK�}�d��	�P	es��/��L��d�We)\5�z�v�ґ��´�c�A��� k���<���~�W�����Ꙏ�f4�9�1]�$}��c���p�ƲT��I��|B�k�YM}�༃"r��ɀҁ�a}�""wc�7H�p�KzQV���9z?��(��joi�΍�sW�f�%,�N����j��O�I��O��������)M?D'��y�c'�ͩ�s*\ Ƹ���>�'?�t���2��H�G�$c� ()p~�N��V��`nc�R'�3��D��$��k�P��^���&&�EJ%��CH5�%�V��ӡ�E��c1Ά�٠���2=���%ÅrdJ�����3���)t\��C�Q���8 ���a�,� X~��^�@v=�
�����f���I{�}��D���o�L�\��P�#f}����9-�EG�c>����� 9ʋD�E׹�nD��3�c׻�
P��j�~�X_��sP�*��!��YU&25aL��r�eD"���~�U���鹯S3�p<���P-w� ���~�������(��Oɇ�k��U��:��C�~%�L�0������2�������N]��<�i-�9��;ya��94%]�.2 ���D���P��r�Ʊ�etN�S��q�Zɮ?�Ez6�����9�
����6��b�'2�_��������+kH���|�5!k��hV�xƧ(Ue����S9��MO�Q2wUYbV�T�2�k[�[���R�90�Ѡ0��P�~-�v�&c?�ߐ:U1<�-�8��*��$W2*ZΌ��9�
��.�k�������w��Y��M& #D�¥,��q_�^e���2c�s?\��4�?`��\$x+h��Ty��/��6�I�"��Y�5w��D]�8И���}���l��Z����}+���Uf9v%�����2ФQ��̔�0��t�:TT�,���h)[������=�y��c�� v�����QM{~�h�KLKoG�P����*ui��T��lU����ʎ'z�]�0��0J��B����Ť����ZǤ(DJy���a���)��RoM�o�w��(gP�U�6W�5bC�ث�XȰY�m��</�ܷ�:�O�z�NS���ې�Y�g�B�QPR-lK�Bi��Z'��z�=�r�3V6���V]���\Ա�C�y��!�fI���kH��>j��o�u�#�4az-	���p)�\�ei����V�5��O'����eȞ�Ъ�������.��	��������d=Lο�x��2��i��/�����	*.�������IJ�\�K	�bD��N(��N_֡��U��!+%=�f�k �m炱����B�0hԠ��Y#,{�]��4�0\ )wx�������^�Ѓ�fZrHx�*S�e�kŞ䰃,�Z�P�s1!mǷ��g�Hر��1�����PL�޺LN��R+A�R�a�� ����s��`��g�����z2���"�-�afy�bh��,�o�h�YZ��b.��]��{����x�1��k��0�3;@�n��FOf到� ��v���W�86jy�I-;�3����~����g8��������8k����+��_9��_�=���Y��|�H5��=;�n�SX�����dGt����i5�@8�Ж�ިX���g}�캈��h�R|����E��J/� y=V���aĮܵ���x�=���y:4?�T��O�����kǎ�[x��Ž1���pw_:�q6	�迓���#��]��ݗf��&��IE����^���B�aMK0D�#K���2�1�k0�ٔ�A_U4sb�U��*6��M%BW����Y�4N�.�	���m�_�b+��q_Ķ\pq|�N�Ǿ菮��z�T�.�	������ݴ&�UO��k�=�_�AEu꿪x��%�P�,s���$�p�y�E��V�0�oe�b�oPm	��v��?Έ��V����^e���:�������%��5���8sC\@�L�\�t·\v�1�|j���>ij)�`>W+���`�k�D��-S\%����M��eC�)���c�x��%���Fn���R,'���a��-�`v�#�3}��3Z\�Gk�e1�a�l����gT����>���q��n�x�

	1��{�3�{�]��9{K��	�@��
���M��O�/L���M���ύl�.E�bS�� �H���9jQKDJ�ne�U_NX�}��2����cc�����r�r1b	X^^.~2��>T���=��ʵ�\����L�ݯo�-T�DˊM��ފ�^i��&���\�Da�'A�$K2u���mֶJ��-12&&��1�7���/e`��?�>�S�e�Q�Y�U�V��%8�_z�1�����U�|T���ux7,���������j�F�WB����E�����OK�������?��?��������g�حm����g2+��8���#(�+1-�H��8>B�B�UB��2�hהPB��3����19�E�;����}E�7>yO�R;w/]�'���K��h���>�\}�v����/ND���(�r�4��R��r�N$C���T �m,|��v���R4L���фM�:�>~�����7ω�4�q��n(.�֣[���պz}���Ob��w�-g٤�c�����Xf��q��J�i������=�!�����tg�;�����A��c�l��y`�]e�R/:`\k"YT�|hX�/B̈́4�����jω���Z���m���&�ض�����[Ô��ݯ���z����ve*�'�w�^,����N,�~�{���AW~���� ������OĖܓ;Q��ЉC�.3�/�+�lj��1�ؖ2<����A%�/����Z�~A|e8�D��LWqZ-�y+���Q��/�1����Au�:_9�3�!9{�b�d����婱�@�lG��n�
��7;r;���Z�IԾGl,3�H��?�!���O�C��Y��Í�oO0hL5m��~T혐�|�5�nT��q�[�����YY��l����O��}�6���t@��O�Z���P o�����g����gr��i��ӟ�n�?���D_/ ���D���zg�Z�idzD�/�u&�/�:?��Ոsē�����hr�,q���y�c���αo�ln����fb�����;�����XqJ�L��?��`4�_�@%�_��������m?�%�
*^
lGh��[�T/��}�_-t-|��x��2ڸ(��Mb���r�����OxiA��s��M�:�G	��ߓ�
:���mL�IO�{�I�?H��tR��
�6Z�G�s�	�Lm2#aY`s^��C�6�i�Gy;����U|��γ��Y$K�����6�j�=��Or~�/�����S���%s�hFOX����c���x� U�����?��g��I1�4g,;�K��#��05�՜)�To�"B{Y��Gzs3j�ú�?��[�6�u�]�Y�9����Ũ�a?���me�]]��94�9܅F-�B_��h\_����G東/_'�i�[�x�)�rn�Mͻ�r�X�2�4�q��%�/�f�y�jH�"�Mz�
J���l������lR��_�=6�茺5i&g�LB*uCg��0�&D�hY�S��l}��VA@��D����>�ͥ@���T~s�}��މ�tx���p���q�!�R�٩7Ʉ��J�7���n�Ն��S�~��8��aR������m֬�b�~&E�����rq�g�C���}u�W�j&j�O�;��D������zr��o��H�(�|������il�;�-��}��w�D�i�X��,���W��mwB�ܜ1�9e��[�^�h��蟏$�k&
g��YD��X�"��q���18�z�@,��▓4�E���܉K��uV�T���N;-f��f��oC��IO��[>�+�a�t����U��iA�D�[E[��jh��ƣ�ԋ,/w�寐BZ����GJ�5z[��>�TR�r�i�U�>6�1E��ǳ��(���כd�:�)'a�J�V��s��jN!	��:{!h`k�x�$
��"U�m�ơh.[V��X����ΚM
:f v�����rS��6���w�-ھ�/[�/jJ.1�GJw6L�R�RUWf�T���6�����X��u��<�����T�9����XB�2�Gٙ��؅Q�U��
$� ��7����@ qY�l��/o%�D�P����X~�Dw��h��w}"(�q�\ջ+n��-HǋhLfxv $?��Й���D����1��Fev���.L̀��A�,�!�����=>,b��AO�Z:c��}�M�^��1+�U�ՙ[�RE��g��ތ�~vS��[��T���7J��l��.���fqȷ�2-*�iRC�{�i�1�������8��<��Д+_�v�E'!�A,���e���ȎL`�J�\���5f�¯����/t1�?�R_+��+"�2�7�s`�ki��}u�.��.��K�b>+e|���&}[�h����V@�א�p՜�	����.x��z����i��&_��\�n =��.Q¯�1�OCe6�}6]l�A����ͨ<�d��1�p���bS��u��	;�kS����������������W�1���mX#'�`�r,����Q!Ĉ	{�W��Ȱ��.�)�$ljz�˗��y��S��l���1{(a|╰f��w����ܛ�3�p���~l(�rK��)��N�l�mձ�K������R�h�3�`��a�����U�rub��0�!�O�+%��}�̊.ݠ��B��[�(�F��(Lz/�n��T��2'���Phk��$ ˽����!�n�ܯ5"Ν�fLpXq$º͙�ax��v��ծ�~�|�V�9òc��'?(��
ԭ̱�*�8N���6l)�=9�B�0>=9�3H�V�R?�z�%�K5s$7΃�I�B�fj���V�N=���L,raAӼ�
�x�a#S��
����q�Hi��Չ���߀p�Kq��#?��vm��LX]���=ej��bi�l�N8l�ϕ}�q|8&|[�?H�Ŧ�G�N=#�A�Y,�OK�u�x��ᤸa*���?�"�mH<�m�s$�)��9�ߑE7�����B�Y��S>��?ĝn�-��A|�O��r�>!�dN�L��?�^�<�t�#m�G~(\�+�E�x<�~.�<{Ǳ)��K��O :?T"}D���p�\��y�q�T�o���ʛ�ג����shu�W�'U�s������5K��<h�}[sL¸T���hB�Z(���N�D��Q���T�N
hξs��s���/��;�&��^�}�Z�a���3̨�o��=�L�
�{ç�*���۱Ŗ<�u�����%�MTM�Z=�g�4�!W�P�)S"z��H�{^ϓg���1,ŚI��'ɩeia���nB�v�-_�<��T;* �}�#�M���͒ח�}�?�Iռn& ��>����4P.4��h��@I�![w��9���^�`��_CD�uޖ�~��70� ��!&�2���k��}!�~�I>C��᛫��gyv�D��I�q����m���[y�ՒϮ.f��5ka9�,%��t���x��(0��C�*+",��=����0CW� "Ӫ��ݮ�����Ge�Y���q|��g�A=\v6݋���N��<cm�RۺN�ٳ��)C�pͺAݞ ���[�V���S��N�!�~����e��_�a����>���z`�WW�+
d�C��!���~����%��� f�VG�(�Wˤ$�/
O�2.f���V��W��}�k�Eԏ���UgD:n@��a��~:���6h�ϯk�GuZ╎��t5�T,Tcy��������Q���m����=k��4��9q�*3�_H��q��c;��٦��,m����(�
�|,s���e�
����2��X8�0H��Ɉ�KHƦd ��jvSVU�G~���CZ��eXE���@U�{ٔԫdP��<��~}
��k�V�釟����d�3�|{��{
��?��x��ti�o�l9��3{����̏���R��vp�,�Cy��#�\��{���6�e&ˇN}�ed�춭t��.��u�6�K�N�4 ^�*fTw���U��u�詚��)�*���<�s�����F5Mҵ�܈ j�-;�h��~	�OR۔T�)'������Q�khL����"#7M�u���Hi�ڹ'c��=+:?��z����U��Po����.)��ʵ3�<�<j;=%�Z���+�P8hFup˼<o*1��$�q�*plUPFZf4M���j�,q ��26�b�+�@�a��[~ئ�c�m�U�R_?tt������c��!LB��9h�D��je.�!����%���-����M�����{��t\��V3�j�S#{�'�v�5G�<�> ��u�%=K'N@�o��^�_��&�9�>҅R���x���B�js�04���O��@qҫ��Ɠ���J����7��Ep����	��HY�\�j��Wq�^��_�����|�ٜEZGvu�^�yڻ=���4���Z��[Ъ�w������D�� e᱊�=%N~)���zji,(�~�N�t.4�G��M4����|�\8�$�VR*�f$9LX���:�4�0���Dn���R~���B{_��̰�� 8Pc������:fͣtU��NUULps��(�|��w�`��[|�!%���~��aA�p
���΋nE��[l t�cU��׹�;��ih+�y�@�����N��[~qPϥeY≰��
�8�Yc�$&�؜�9�kj�2�K�O�SP?���T��C��'P;�sD�1G�n�QiIr+�cU.�B.,'���uU����nb�\\Z*r�� �Oi���
h��0[���Pă���WI)����F�4`�n���L��Oƿ}�t#!ͧц��}l!����Ufc����^m_��Q�����@���� D[�N����#A4M�-RO�Y��7`yO��D��(���6�-�F���HbR��|b����
��+��g �,K��:8p}����7?��0��]˩MGa&cu��Ft(�j�䇞������qL�ӝ�t�ya���d��V�`lh����Vg/=�́��$(���= ���2X�k�o�)P6��ޠ�7i�-�+>�ϧ��a��o�.�����Y�i�����R�U�Olŵ�N@�kG���0Az�^(����XE���?��zS~+v*�j()&e�(�A�����nn!�>��j*)0#�s������a7�x� ������̉����[��eC�I�xq�T-SIY�崩c������;fR����sm>۔H_zo��_`u@_D������Ƣyކ6�QfH��޸��TS��|#띺ܹjt[~�o�Y�R
�Nu
a�Tj�� ����K.q�w�&��粼(��p�N��O'� ��Le�'˾ڔ���eϦe[��������#ݓ��Y�t�UieP�t~�'_�B�B�S������	x}z��)�U�8i�Nd(h΀
1������sQ3U/��"ʽ�L^�d�7�K��(����˄���&#�� 7��m�g=ס6��^*����`>��
��V�9�̷���&/ٿ�![��[��w�!:	���t��ƚi5I\4�E�9����d�n���$�'�ʗ:Y�bퟺ1�l��5�y��ħl���˻4�JW!UNZm�mu�?�� �(�JV�Rp8�#'\
��,�6��Hf�SF���x��]Cg�����R��*hIjK�Z�̰N�W�@�I�z̷�H�b�⍟�V	+Q�-�e/��U��g�������;�H'��e^ӱa� �i uK�_�~�B�H�y4��{�y��� ?�q./�u�_[e#�R�#`:�E�|�a+�~^�R�@4���� �D�=:�WPc�Ҕ���ضP�y�TA��n�h�S���a�qu�t˝�*m7��N�\:䷥d���+J�C�Pa�*\I:tM��.9�y��r��ko��	iG�^�7�w�N"�ԏ����}f��j�Y,4Pz�3`��A/��m�
����ގ�� ubL摫OK�q�dq�J�CT�/$玲����Mb�g���
͡�YR��/���/mTd`7�n��d��xP�)Q�W���ؐ�wo�����9ض�\ ���wS�:Xji%ᤲ�X��-C��wÌ�:�e��U(߁����%�?��#�y�iׅB�� G�Β��|�`��T�TGR2�{��j�-���`�h����:��ȧ�.���C������P�˗�׍���}�~��xt|l�Y�9���c�!L�cIs�Ҳ0�;�[��2���4��������gQ�����s��1G���D��>MR��۱9LS��`����f�|���	�Lʓ�UG;��;@�q^�4����w�|��+I�.�Ѧ`'�ZͰ�g���$@,PXn#�-��蠖H��	b�:�[H�}��^���pQ6��������G9�w�*�`{3yh��^+�8)����l�.����/�a)\�]�*�1���'��h�i�A�SM�X� �vt�@�%�k)fa�Fux�kt"1?1�u��pV��Η'���Ql{�Vڷ6^�&�B�[����g����+�F��}w'���	e��*�~ЌY�5������z�Wf1�uy�E��s���?��6���XB:���  �uA+���7�����+G�T��a�J�+69��y���!*�ѽ���I�J�Of�a(�\"�͡�&q��F�p��>}�jf�H���|�18U��DfbOl���1�(A�H�����V69�G�����k9���?�mh3����~�� �R�zM��	� x�k ����@����GuѺO�D2t��m�8k�t��mщT�Ԏ,�p����5ӎ�<�mX�ba��6tT`��J$r�v7M�(��m����"�:�����u�a�2��{�tSt�|"6����EM���9�-s�3��lE�+����P�],��=��@�%��e0Q:�~gށVtr�i_�IKmQ�̪�C���OȌ6"o������X�uF�zeB\N��G�D#�c�V�|�S�C��m�'��P�'���7��u�C�2T]�)�~yX�R��ab�x#A�Y�؄�����Ne���Z�.����8��?М~�m�8�?���:�їc\�r���\V
�إ��	�5�^���m\v÷#4�_	�Eԍ5	�Z`i9�G�Q�I����t�o��d\�i�
k�C�����b��M�iuI7@���8?�*g)�<u�����6�p��G���<=�� 4xg�ywM5��%7��4ԋ�1�(���)tnO%8�d���d�l`<�d�4��!�;"-e^bh�:W�s��۔3�h�e.�L���������!��LN�*u_r�oR#����z�9  �(��r����<���Dv"��)k���~ꑺ6����PE;�Qr����q��L!�ۏ���Ay���H��A_�)��&�l��w����I�M'���PQ��f��\�XN@o[��<�
��.����"JіD����bX��:�`}�n�+����.wծ����"I��m�0��®pZ`�u'�8ծ�i%1�+�[�'�@-C�Z�����e<�T8�1E����X�����]��u�4�P"�!M��k�����{�n�]f�	��ֱn��ׯ�Y��"�*�>���6Ƈ��D >x:�tbLї&����A�8>���gh��vf$�j�����itYQ�ϙC꼶�F?�zkZu�r��Nӳak��k��,����d����v�h�"���{u��bϽ��������Q���!�����Yi�)����~�l(�ӛP�[�"��[lr�Cy/�F�+ؤ��6�sJ���;vN�Ilz�ne����U����[�	�[V��)��#�ޛ�ei}NQ���B���\"m}zNw���`�Ƥˢ��ո����>{w�/�� �,�J��]����C6vLUp�p��A�z��ą����^[T]F���ͣ�S�M7J+��T
+3������p���u�t[	���|agjG�|Lh��{С��xoa]��"�J�Do������;9�<۽]󳶞�Kȡ;;���.��z�ۄm������UO�DR���[_p��\��Z��љ�3c�*S>�XyjtU�É�Z!��|sɃЯ��<�1#����L%�Q���Ȧ�iR<�@n��uwJ���V��t7�dt}�v'�(u���3���;ەߘ���LUn1宧�����26����W��Q��"�s2���x�׈�	qƽ���e\������7������l���;}T���,L�_���ᰲՊv�<���u��u���JHZ���S�Q������."�]�FK}Ɯ���P�C�%��35�V��#�(Ƕ�ve��ں����%j�T��o�������\�C���$Of���=�2Bݠ���PO#)�z8i���D������X��Z�&$c�������V�����6�,옍�0��U
8�57ֳ��?��N�� +�-��	��4��R��l����`�/(�mU��6/"	d~�ݾ%��rw�왱6@ҫ���L-���B�͔�jM�F��ׄ�˼�ݎ�'��]{IR�5�xam�Ys�4���͢j���3H2� S�6���p��[n�J�B���sl{`�6�9r�J�-11��EҚ/\\q�1�u���C?{��pS
�xr��7_-����dn.	Ҙ���U�8/�:�l'��d��U�Fw�er��J���?��يl��P&}b	��YX%i���fz�,�������.������Y3�sU�%�>�j7��Hh5W~'6�)��Kuh
�N&�����{/M������C�2�"����PE#��=i(����b�d��W�Z��/kG���
�9+9�a���H/�����*Z@d�즐�v╽�PDy��/�a��5s���m7(&)�!SAz��wy/_����{g�=�	\X��e5�xA~�Qw�S�����O��p��`�����B#oV�V��R-����(3�읜��EE�{+�z��Ā|��k]WT.��ӧ��k,ct@b~���g�WPA���m��/ވ�����Z�T����mb�h�lx��3�:��*v���6"�s&
�bǆ�C��Y����f��}��F(�v��v���{����,�������|�SKcoίz_o"G>I���5��хNc�Cw��0	�bAm՟_�����$h�[Fr��{�MB�i�oVlͷ#,p��w#�h,���<c���H���x��M�}���]~�z~�e��>�@��;�>&3�k�u��T*f�bt�^�#�xv��b����bE~z<�O�©e��"���Y[oM�F~��˸�j2VY��N�bMx��l�Wmkh�Dm���p���� ��!��{a4僥}� g��Pg��j��)^�b32�a��w�t��M�03q',HLL	H�\[b:�h(��zR\���;}LS1�b�Cp�U��\Ut�bݤ�B��EU��:͖�kQ������5�e
����?`���S����8(�<BV����C���ǝ�z�d�5���&_��	�t|4�łH���f�Ά&^��k���U"~� Շ���X�ʅc��i���Z���i��Z�R�\�f�g�]�>��O�~0hEsg�ě\ߦ��S��Z����A�]fD��h��������o�����d|ǔT1���H�7p���b^����_���$��SS�$;��,���v��ɤ��G/s�=;��t���,�<zVP>=�J��Z~������1{�yܻ�4�VyGւ�|"�J��lqo�� ���.��Ü'�Տ�ֹ����]�h�i�������4{�Dp8�Z�<]b���.{y��1j�����F(��T4O�d�3u���s���%w/��L��ֳ����[u�\x�����m��*���C�pYp4��gB��](�B�?�t��C�y5%6���0��чt���a����db�QgT<F-�쮍58ii[�&����o��H?;ĪE$����TX�73����l��ɴ�W�V쁪�����O�|����:�6j#�V����4�Q��9�{�j%S��Vl܉=�(��j_|�x�VO�P�G�feK�_MGy�q\��3o�.���"����Q[��j+q�W���ZU�S�	�^��M�"ի��{�T�c�3��������	sKn��%�BP����+{.�	��4�ύD�L�<���CΕ`x��^����Jr�};��reIƄwO@��{6�v�R�G���-��>���*6#��u�c�=��c {�̈Ǎ=���}u��Խ�z�����tͭy���t�׌�ߒ{�T����,��kW�����T���C�aIIg�Z��s�$[X�b��tv*+�qB"M<ͯ����V,�OTfK~ݻޟ��z��N�ŊE�CJpe��(�̱�/HL�O������O'�[/.��҆���+h���nqOav�#a��rۍo�zgg�MMz<Ή������e�(w���4���UT$�Z9�nʾ�C�Gk��:*vRC�/��n�?aR=���>s�����1pS������ݕ��<�g������;	�rm��%,���K*	���J��mX*�w�Rǂ^�q�����R޸�{�<EH�H�����7�[s;Kh�tW�?q�O��C��'G�W���Sy�t�k�z>lq�A����Yk����,�]�)�\�1��D���z4�%N�$���m�m�$�A���x<8��m�Ɍ�ʔ	14�i�3���?��pp+w��碌@��X��t��\�{$��Q���wf���obΥJ�=Z�z�)�!�d���ѶB3C9��g�#ḡog��cd_S>��'��w���n��dvv� C�m��%=@���R5X%�ٕ����=9�E�ШV(��=�� ����+g�Sc�b��+��.���-a�x{y��.��ɟ�:��Qm�'r�#5=+�V��l�H�(���@�ѮԨ%��m�b���ߥf��W	䳦W64
eu,��Us�7/rsSc�WGƍ�����,8_4.�p��G�%҆��~��9��6>��,R %`���]N�V�F��HA`��Q�8��~s���ߝk۵�Ru��A��k���q1N����5ImX$hv\��uD��ԑV�_�2a�ۺ�I�Iw�32���L���x3��H6��������2ȣ[c���~ye���`Hp7󺣜q- =Ȓ9>s�zH�t6~&E˹.�%��Ҩ/c�U�E5V^D�a��u���N�K�7�Y������3�w9þ��ߔ�u���C���2w�c���]�fK�J��Dk�oV���n�i��v����g�I�춳��H[����<����2h��>����*_��r!��˜=�}��k���?�Lx>?r1w�A=�*f�]�i��+���?��Z�j-=�[��6[K�s�ۿ�'*$�{��J4���T�Hx�i��写��v;xs�G��3P�9l����+��C!���^G+�y��Q��!�2yZj0�M{��$�==Á� ��߁�T�&���|��kC����'��S����Tڸ��"^zjB��@��i�u u�$En5U���� "Pu2-o=��������g�j��M��*[�6���l`�Qj� �Cc��^��/�昑(�v��S�d2Q�U�wa���ϿjP�i�`��HÇ֍j��Q�G��fY�zZ�R�(-3��8�xX���tQ��B��k�{�U%�iq�7z��Bh��g
���o������k= �u�Qc��S��4�� �c�0AN�5W�� Yz5�g�T5h$���h4bq�d���1Z��%z��i.c�:�uC&���Dzz$�E�`�߾g���4�?�l��w�]�o�@���/fkeU�{�yL��['G�5`ԅBCӞ3�8a��,W��9�$0�W^	|3���E�7���8ػmX�����[��ڰ��'��e@@ ������3�,gf�dV[k�HQq���y��� �[g�A�l�XU����6�:��_�Pb�3��k�g��[���D��p��o�NlPU<ن��](;g̾a�g`<Ei,q��?c�� Y�م�V�@^e
Xy��Z* WZT�4�[�!~����O S({�po2�}��bD0��J��CO��Ae�laV�"�so�JBl��U"�%��b�-+�6%�/��j�\d�ӳ���t��3�����_����D��� �Yx�0˝��]	�R���m��R���᠒-��������w���V��yk��-o���Ox���ڊ��a��QU�E�'��oC(��v����RjB�v�?���#��x'�Wa�\mљ���e ,W1X�Y.彏�Y��I�f��XE��͞�tW��RgU]
*���|o����w��N��j�g�-�H�:���'���=�_W�MX�i��sת�ً1VQ\c).��K���[��rwm��_\�k�[D����$~}�������H}�3+�K't>�O��a=l������.=UyA�	Ya��tSt�R��Y�;W���[4�&ZՠǛ��)�	���cr�@ݻ?ݑ���ͯiX����$���=Y
���^�q�]c�����>7v�����y�Q�J7�E������?S�-�^���B���]�M,m+��F�+A��[�].N����ȯwIow|(�Di��@Ttt��ґ����:�+��=P�L$�H'�!����莧h��A^�۩�yս���/횑S�w�Q�R��bc Nʘ�3���P�j�rϒ"��X��R���?�s�h
Ι�Ӯ���[}�;)����5@���6�m��2�$����r�������z��Ǳ@���.E�Ai�IEB	)I�R�F:d��iF:��r�{�{��������7�f-����>{��y�9 �-�Ij�_����a� Z�f�4͉����[#�7��P;���;��:s,R���X���l V������~O��߷�����x.�l�&��9�����=;���JBݟ�7�V]�MD�Ql�ت�Ab`�̭-�7M�R��E�e�?.��v������`��\%��$iq�&h�|0��a��u�g�ڨ��9��T4���aK��`�����cqNx{U��[�ۚ>����?���&[1zQ�����h��A��I�V����D<b��_ ���e�� �1:�_���Z/&�)�u��2�!��������{��b���,&99��'��쭿{V:Ŭd���G��z�g�P�8������b��	�8Ku����q�Q�fc�ȉVq`�7�Ȫ^�>�4a�IV��l9��ut�B��Q��v(_��q���ܼAn^`'N�S��4��4��-����ku9�Ȳ�����S�p&1��*V�����J�V�Pkh�㟡��n��hۼ*e
��#_��UW��a*����3�0�еd��"�c�q�?"��Ā�6��x�:�3���'�q��A����X�ٕ��y�Zt[�hQX`7�[��nC\S�2��ە���N?��+Z!ۊ;$$@(�w�}�`R�X�Qj�;��=(�=:v��(�Q#FGk�a(�sjx��֢������HL65�I�-j5��N���̠�%J,����ϛ6r���ѡ�%^H�6�Mq�޼���1��6���H{Nɖ@U`��"���NL&|��2{�Y����G=�c�!^�S�F�<��(*�[re🡶���,��Q�����p}u�ͳ��N
�w�~|�ڋn�j���,�j�Np�*�S��o�KY��fS���u�T6�#w��wvܷ�I��ȑ�i(��Z�<�0�'��7l^M����]]�'�z2�O9h���\��0�k#d�R������fqUR�,j����ΆoT>���I�D�ƒAm4f��$�V9)��f�j�=��A�vo�Ǘ���O���5�Z��<�\¤�&z���/F��V��h��9��	�Ye��Q7,h�VreG��  2Z⇇�
q�_�
n����#��gf���'�P���hB@㝂�Ҟ��ő�X��Mݡ*�7v{�l����dY����WQ/����ɓ	V�����"�r����w]�O���;�J���v�L].������կ�2c���X
L�ťƄ���5���u謪��@��|0��B����?�T���7��
8��#����^`}�شN�8�a��'�����B���'#E�/vuJ~���+޼���hމ�IIv������e	U๕����a�ǍU�A�#L�&j���,:�<]#Z�HB��>_���y"/����m?M�I݉s�W�d�&Z�	EA�1��^�w�[d�w/m:�o'��Jl�G��o ��T�0ub2U�ٌ�6���B�P���Pm��T��H>�����i�`�SB7�"f1��M��,b�U�+�_�\G*Z'K:Sse=�0�S��l��˸V��5:���r���C%�+������hV�iND݆Dw�K��t�C=TU�E�(�!}�8�k��@[M�=��"��"���Z��T�dr���_9̿�C)ƫ	�5�9�����x�����ɻ�gs�%��!`�IN��9 <0x�~����s�oŏuD�Bύ��:����������.%��G��K���E���=]�0�b��FU\M����dj�7�qo�I�46l��z{vVr�m�jBC��؞Í�;��h�y��̔Dv�4��L��x�wc�V����d�0dX��z� �&��s	0��{~w� +]���Ҷ��������Sd���Yԯ�����E�>o­	-���K c�}� xd �V��'L������ŷj5X�������q�yk�TV���7����=K��X�L����p�U�D��P��g�~>��8��M�q���q��?GM�$5'�?��7�?'Qd�s���Γ<!��9����9��q�������~��E�9*"�y4��y^�9��X�o�>F.֭�nӛW�p#~m=�Ճ�5ޭ�m$��ͦ|�fX*�����P
b���Q�E>��)׈7VJ|�O֟5r �R�DY-���ah�6$�V��\�9�^��0X��,!/�� [� �I�nl�t���b	@f�����*m�s
JPP�xOO�xl��@fQ�G �̻Uo9�GrN5"_��P]!�G�,�;xhKU�z0kE���*/�-��]� �Sw�^��������q�����S?���+:	�[Q[���%mL����'ۛ��W7���lp����b�_!��i��H�U_�/�1\pX91�� ��̻�����o�'�ȴ�%[Ͳ�jy\<w*9��i��릦��P��?x����()�����A�A8[��}ۨ�P�=���xf'����.���>f� �0�,�Q&�����3��`�'02z.'�b["	�q7g��&o}�sV�Z�J�JW�Qb�*:��A/�����[K���:��n���vf�sദ��q���m�&yfQ�'��/{"��_ϻQ��#�d�'�.�ʘ;��)I�|�q�8���jG��A�2C�6�xz�Ǭn�/6���Tq��l��~Y,
���`p���s<|Y��4��/��p��Q\_�9�ԠJ��~�:Ҙ"�ԗZW�����\��Rn�M?�j\f�N��@��5�i�w���hw�C\���!���rM����,9��b�>c�S���O	h���m�7tWY�΅��T���0pH��	��b�s�mA���շ�|$K���A}����R.��uK�ʀc0�J����*��
i��t4Eq�� `�4�*����kc�X��T9MM���2��w|�����6���ۨ�4��l�(E|��|�Q�p��w��ab��ˆ[o��*9iͶEg�[u��>3!�'a���T���D}� �����āo�5ޫe��:f3�\H	��?QD�ɸ���Ccկ{��<M������� ��T�n0nBh�"��~	�~gc��Т����}]��NS�C9q�����[����Bڂ�������ӛ����	dS�Nv�c�ĉ�3ZƑ����<�tt�B���f�X��=������������Nb�Y�Flt�J=0�+w��#@�h}ON���I��i�A�.N����x�|�*sT�`�i]M]*�@ᚻaú:�Ƌ赡���ޢ��b���e`��> U1yN1�	QL��}��?���<8@��J.7 ُ�r�hH�P�����H�\�͈́Q��o�xbF/ب�����>��g�=��o�mfM#Y\�n��>� �!�ie��K7�5F�߄�cJ1�K1+����9����xZ���.I$uJO-]�b�ȮȠ��ǘc�!v�3uV��4nJ������'�[Op=Z�Ԋ���(��waD��{����/�W��MN^��jQ]����}5_`���Qf��\�1�}�̼Zc�ևM��s�M5��|��ߢ�B��4�1�{L�4eE:�TT�(r�h^�KQ�0���0���F�m����l�����|z.�m�Kʞl�_��]�_��r�T�.{��H�kq��u���07�b6%�(@(��C��%��kO�R#J�}�;�67��a|���1;���)�#��&�l��6�߽�\1+�$&'{�Q�T?/c��`.�� ��"aM�2�,E��ĸ@4/��(���0��UYcn)/�f�������,�'�&��~~�{ɫ�ǹ����Z���FO�*�����􌾭��[�zs�N[�4u/<��wG$�ߗ81�9`���gh�j�Z"��i*��� �M�ʁg"��\MF�9!�N�HG	 �d�m����Q穡�'�]b������4� ��|����髟���Ft��$��
>��S'��[+�JI$�a�v�����U2���k�����nn~�KU+���I� H���h(y_`vO�� P�ؕ��V�.؄R�5<(1B��@������0��t� f�?�?�݊�r��@?����ZIh\
�$T�h�ߛ��)Q UX���)�E������T�1(���͍#U]�)t������`@$�z32��1k8�c��Gzq�Kߣ�0��b��#���ƹZ�>o9w]ii�F��8$ܞ���<�)q����5)']�y�u=A\7~�t�6[#�,�Q��v���u('A�s+)~�&j�Z@����=̇ޅ�'vtts6�шNC��Z�b�9��zu�G6��|W�f�z�hN��^ڐ�O��e�F�s97�gH%��:�?���Ǌ�i�V�TW�`��"Z�:��c�r�A�v4��,߁~�i�<�-g����lo�x���0��-:ij,��3n���#�/�G1���DPK�� K+������p0���>��a���f���^���/K��yR�
�z�2PLJ7k���2�\�MY�ԧ�1�G50��U�{����4Z���V�M/�;��&V��J��M��gݤ�S�l�t�s�xeL�C�Y>m礴;:�����fͥ3����� d��9}��w�7��坼�b]ыm����y����.V��V�&oϗru&���]��"r�w��=�gR������;���}ȃϬ�~w}��7 [$niOK-�Sբ��4ɻ1zG��]�b��7x�Ž�y��L�����G�����01S4kg���Y��/��q�N���?� 8dx+��^��-�{<���n�����oeaF�6��ۍ�7�����-Ƈ��}|?��\����n�ږ�h�YJ��x��B|$�~�ҵ�uMT��8Bީ�<���57�^yQX!jI5��pIx�j77����_�0�&��FM�XS팧,uC�:;��Lm#=��ބ"fS����s *�@aˠ���w����u_'h1�=q	sDA���� m�k}�_�pÝE�t�#��j601�F&�(I�~. ��g�9���e���z9�8�ٷ@�h'��S�	W�2�ă/e���D�%i^�����o��%K1�����?�b�� ���� Zuy�~�Ƽ>zv�=�'؎��;O������K�u�������]�p̐��z,�ѓ>�	7`Wn��b�ЧML��*���\��'���A/-N��}�	mx��V�6�)�K��ŃEr�&��l&�K���J������~��3fE󘕔x�^zT�E�-�AO�ߓ~FC?^�\R�H�����|UOr���~T�3�h��6�+�jxѽ�U�����@��8�B��6�,��3�Ɵ��v��H��xn'�JB�O�'�Ę��9%�p�����m�����#j����a��I��Q�@�
�t�[�Q��J�B�V`�Tc:i�H�k����Ȋ�Ut�]�6w��fP�6(L%x��"[��.�nxOꙡ��x�L)#z_��J@z�"��o3����y�N|=4����6#�-Y1h���-Ɖ�����S����y�$U��N8Յwd�w�����Wt!��d��7X������85���TrȦ�SC�OFurw�\/���º��j��䐊e@I]w^b�L`�J5:,b{KE�w�5��Ou���=�Ŀ�hױ[��q~)N[H���$��&mD{����'L�ml��>#�-ٝ��T�-s��&�imhV��/q���y6U���P&If�-W��y����1+�c�"��v��͇'o[<�Q�D��j X�n.�ޫ���;j���R�y\�������bo͡i<�㙙�5D�IfUý������_{��g&�8�OܺǱ����8�֣0*�m�1 �<��M6Hn{��mm�h�S�ng���3�M�臚%�MSP�y,��JV���a�kEl�E��R�s�NZ�	,��U�Tr���:e'lЉ��9Q��%
6�r����AuT_>Z��y�SmX+�k�H�#�ٗ'�t�PB��kr���9����MGG����w�f�~�����������g�'��8��x؍'l2�S�ѭ�1N�9q��輮��6���<����N��R�鈴�貨�[$��1<q���If_2�d ��z��l�I_���r�
bw��;|8�^�����m^{�
�MI|譮���tmM==+��� ���J�n]��F�Zy�ƥy@:1Mr����v)���<�ml�D��љM��^��5����B�[}�\#��,��������S�^5L6=�)�
'�ɜ'm*&\1|��ik4&�ְ;s
Us�{�������sM.TN4�?p3���>ps��vm�F�����ܓ���ֻ�X����h�(z���r�q��r?�-h:���u����e�r�h�'{�x��W�b�5bD?x�yvݕ���7����6���r��r�C�w�
} �<
�}��M�3���r{�����~�i���T��D��5�5Y��(�·ר���Ȉ���H��8�V��Ό����"T��Dc�1���2�M\B~�:��Wkir2@���zz� �^Ao���m��D�;�qX2�� ���1U[cw#��;χ��:8C�9Fl[�7t��	�N@��Z� �ߒ��y<c-�l��%��5cR�#�L���'�`��9-���8�	��

A�D�X?�9���o��z"�H��v�Y��;�r1T)����x�s������ϻ¯�c�����3�qF'����֦ㄪ	x����Hp����n�]KTo{�`��h�|Tdj�}"��|6@9;H|����r2���9�F�����5������w�����1�~� 8���~�!�Δ��h��9۽�+rz�������~���Kѽ�G���s,�e�Q@,gݝc˵̯�u0yQ �j)ʺ�mZ��3����Mg�o9����+1����O��C�����H��i쬌�,����Ha�.6i���M����W���Q
��) /']1uC�^�v:�狜����R�6L�/}5��V�걠K̩�`Ô�	�C�|�����fy�6!?��zjV���oe&���އQߋ�G�g�1�@Ϩ��[S�Lʡ�ۑf��p��V��@�b�)�RQ�fY/gn�I�[�^�c]�o��Ɉ@9�"߳^���SQT`�@��͏'-Z\�����Na�&�iV�d�t:�<�X�O���:����z�܎�c�7#e��(��D�Z�7]�^E!�(U%�k�]�����^�2k���L��݂J�~���d�N�&e4߼��e���	d��&z*�,�.;��;���K	�v��T��H� A�_���Y��m~�S����%ߢ\�w1=׫���9[P�0����_F�;�;�¯���V�fsY8hޕK_W�N��iy8����iEl���m#�	cgg`A����"���(߲��[>��~P���$����5Z��x�rDn�:�$�O#pz\�͞�=^�'v"P �,��W�?��Ǵ�o����Ы�xٕd�w���vn�?K��nc,K~�U��9˸���Ǵy��(�
2�W���:a���ɉD���^��k�?�r��Z��A����>�fi�������f�װ%���@.3���հ�[�)����:�>7LX��!�Wy�h����Ф�����WG�܋�� �g��l���|ܿل�I��|��������%���|�e�9��җ[N&�܂�	馻C�<@S�(^�y5�+2Pe/3ԟ�3�"��B��Sˤ&KȞX�cz\_����N>���p�Q��ɞ\sӮd6��6���-�/S
�4�2A~�v�_����*L��{�pT)%r���c �Է_�x(d�����a�لQ����Ozuub�9w���L����,iz=U	��Ͷ��x�B��08
���Ezs�s�����q=|�/�T�� O@��`t�"�y1����x��iqJ��Go�pz#�|��y8F~�JE�X�j��|�S��x{	���M����R�Q�<�f��9p���NS��J:FڻKKo����궏�D<g�{�ތZh�i�����ܐMZ�[�b�bmI����6��q����!7��k��n�߹��Pr����3-NvswX<�V�������V_�~�g�U�r����-��/W��S�`�M%y��}YnL���-��J��Ř93g�����"��89��B�I|�]\���Ʃ:�C|��D=VǍ�T���D�������7�2�j�$���ظ�$�:m��?z��#�.���~�B�gyު�Hh���=`{>��;�w�}��p..�����������i�������G�Q'٢�t�W�Х��>����Ŝ��ϋM�����'cD�'�SI�W&�]��p�f/��������iEw�a�?|��!�i4̞xkg%�2[p�aC�9f!�i��m��`*}��BQȂ�ݸ����
��~�B�e�YCD%�o����={V��E�2C�QuW�y��s�$������ٛX���G��^K=sȟw��⬝�Vf�Qo}Tc�x���ˏޕ��[�ߥ��%�?��~F&�>O��9I��U�HYVo1�Y�z�_|:���'T饕U߱���ϱ�&��|�v!�(/�G鏦IG��ŉ���u��m���zu\�~�{Ѡ��Q���ǯڍ}HBY	�����Q,�N�#6�G��L����C�<�����k�Rͣ� �ȭ��	9��1�r�i�G� ���-63�5�BBiB��ת�5G��^�"	�c�ܸ�~��C�k��.�^��U4�c�A���f���� v�d�(cw�ۢ��v�V��᠑���4O I����r4���2%&��%|*�?�MqΊ|���y8�G�]_`��K�K꿎��w�@�vN���]�Y��R�����hoa���YV?�T=�K�>/$�/Ù��ɔ��v@	�j�Ps�㙙�W_w~��B5!`o�U�����ʆ[�W��l��'>�3�K�D>N������sD��oUi�L,�����a���Kۿf�p�P(�dW�|S���AV4��ŀ�pV���Z��fO����H��E���J�v?m��^0�M6"�"T��*��6��%�$ �H�?�$���h[��,c�(�i8O%)^���͸�gXE��8�v@UGy-�~�V�y���&7�4�-U�����r$c�=�����?n�\)ɗ�<y�G5�ZI��c��[��0g���n�����r�z�H����(I�5��+F6�����fL�{�6��ȥ3;�&���S|9u�n2�Yy[]�y)I��1�F�O�7�o��O�t�&q���_���T��� �m�5֭�t�f��u��ȳ�?J��b��%9����CՋ�#���F��d�O 7z��~��3l&H�%��L,��̈�{^ȿ��s}KZ����һ㏃�c�e�-��&!}�W�'	�[�}I�u�>ú2i�=S��Y��:,my�=-�V�c�d�&��%�BT^����.���<1~@>�0��7�V�S�[`���vQ���.x0��g"B����#�)��
������T?-�*�?w�ut��L�Q�6ʕ'OԾ��|myjg;�vv^!U�h���nr��x��_���է�V�
�����N�o�d�G�e���O���9IdW�+}�rsT���M��q�
�yY^�Y��n�ˏ�ik�_|�-������JZ�z��×x�{���R�E���\%؉7���0�҄%c
�&�Mby��3];��O���XX��_�k�3��C�_�o��Ng��K�/q��d���yDr�r�P�w�MR�{�+���w�y/ݹ}r�O��js}��[�����eޠ+�vB(���Gx&|V^8�dX�T�P'�E�����M�0�Z�
�U¼uN���� �&w���M�$-�{K�z�[��iiߘ��Sr.����{�p�]؅�[ͽ��%1ߊ�ӱ!|��r:3�T������d{c�1�-yY���6��EQ�L�S�(O��h�]e��P	T��׶��ӛ��*�ʾ.+��#�t���`U�����F��[̯�Y`��5$�����~�E�{�ho~ >9�Rs�P� ��X
k�m�����DSv!��~I&�
	?���eܥ��Q���;���ƥk���VĪ;L���!q�������E�gV"Y�>�>\؝�+A7�m��c�(r���N���
7��!���%\.�<(�R����r �A,�*��C<�ϣf2䈙�,gf���r�[�IJ:HnT)Ʌ{��E�D �Ő��27>"X�j�6yYN�y!�@W��Ȗ����#ܕ$�(}�6O��e^�rԞ�z��^�D�c4�:L�t��� \�l]5n5�>E�o�iB�p7^��&��&�u�êby��ѓt�� �ͣW��# �����ȷmM�+jI�Q�(C�>+�lgf���u�f��(*KsR�_^yA}j��;��}}k��u����$jB'r̔�g��|[A�J�9�6�?�؍��*b�.���1���$��$<����2�i�ՒS�d���rN\�Nugi��'[���wށk�S��tzu{ �m���/�k��>�d�\��^��!=�൵�`��'���d��Z]Y�_�Ժ�[o��}5�S��#�)����H��`��8`c*4b��|����1�}{��].��Z���#��퐪��)1��z�?Vױf�K�|D`�K9�V:6��Df��o���}�b��6��5S�ȅ�~�s�Wb�$���q�¨�BSS�����W\����X�;��[��wX�Ωuo���8�a�¬G�;�A����d�v]2��9Ju�)�~�A?�b��S�6+�RqH�5���
��Q�>�
|6Z�Å��
�z���	òq�>"�w��0�p����:O�Q�R�/�ll�nG1\q�c{6�U�&��1���V�%{�q�L��y�5*��&�G��y�,��Z�M���C¾,C����~#�`m�[�C��߃c�[�V��i|k�m���y:�j��v7�i����gI^Je�(	n&,)X6����<�o��Fy�;�$�NNO��΍r>rt5ͩ%�V�T�|��=�4��d���C�{�O�����0�]��O���Aa���8�_���H�Kl������ֆC�_��R"�R\��p@���3=���N���I$S�s'�.����2�/ ����L_�>�1
(6�w�;TH؝�=6}��<'�Ē��rT mj˾F�:��[a�)k�3j_XVM2{ؔ���-{^Ha�LL{�fΖ�Ő ��U##���ѝcr�O�p)��g#�<�=�"d�������{�?�ǹ$^ύ�l��~E�G�����mm�����?#킛�AFePH8r�f�f�-wG��[xM1�̅�x����<!�d�;��%����v�H��麪�	.����C�bD�L�ԧ֋k��b���5g�2;{w�A�
ۚ9yy�&&&'�kk��i���}��P'߼�w馟�O�z}Np}��i {�����AZS����|�SW%�h��x�˗��<����{6:���nsb�5�JvT��Ųq+[a���$�L<��'
�V��W_	mI�oZ���d�\���^�9p�����#��?�I����u�2T�Q}*�!aU���y��������G���/�w�F���a�U���[��_<��6���u�m^>������ޜ�|)�>��Ҥ��Ȍ���_�g1<]K�)�A�����}�Bdy2�GYYY�a�Q
x���������ce��gB���K�����=b	�).��5�z���(�2V3-���s��\���P����ڿuv�k�h��M����q�-)���8��!��a�O� ���ͪ58 m�� ɶ�u=p�4��vnu���~�G|�"�<�?�T@�'!��݈��5SE�S�2�&��K�����Oe��H��/Ï���캹�z�/Z"�4�_����L2NEE�������G~��{o����k�-4ב�a�-,���j�T/�0X�D+�W��O6�=x��[Yt-�
JH�2/5!��٘i��sޖ�aV�`b��O�����K!��d hn��ş�
��%�%�V8D���;��F|N���p����Uc��_�Fy��9	v]5@������m�w���#�N�u�*I?�SܷY�$+H��Þ7(>te:d@�;��x��A��M⼐�T�'�j�r�0�E�.#i�΂���O��)��F��xٞ#�~�N�H�_m�${R%h����^��=���g j�a�a�4�؅��bHc��{�ۧ�f��ك&��� �χFF�ǌi�nc��"��Ӂo&+_�����Ud�G�Pg�c�dg^X��9d0�Z�=Kkg�;�߻|A��Ҩp����'G��@���w��RU�lWU �Aȳ�S���`�;,�X��[7�m4��'���w7=�/
�7iP��5�R1��-O�V����w"Ք��S�nM�?S�K=�?�!-T�*�#�\�S=�wf���^F�9]���|T���k!|Oy�f�����[�暽p�N���[:�\��%3��i�8��$�-)^Jp1)�N��C�����y�=�b� ��6HY(C�z辶�5��}Ն���p��7��0V뎹GN���xn�D��3�^H�٦�m���f��z���.Ei6�}���'"�
AYO��W�p��Ԫ+���������v��K7Kn��*���_�£ׯ�'�L�5��gv���Y�$����P��P���Y}���w�z>�7	�Zm�Ql�n��D������@��m��yQ1$)r�	��iS�m���9� do�f�5��/V����chȊ��w�Ą8��}.����@�������6����-�4�)�eh8�� ����}�'.q|��]em�Y�T��k�5�'-�ؕ=Hf�ȕ�3j�R��_�/g�딾�J6��#I�}�@��d����p�y�K�wq}������j�g1��k����A$b��$��0D��ȈVye�|O�e, ��6ާT(�7�L���������2$2�����W�? �8*n�
}�u�@�%���'��b�����H�j��G<�
�J�������o�D���r��1�z	��x��,�(+ߐ��;�`{����t���a�s����g1�c�+7��;w��WH����ݮ�A���A��𮡜�h�[0��		x>�5�f��v�K�D���~�g���d kw�o�
�Y��wܬ���m�}Z�)���+-�X۴i�>��G�z�/'5$��E�v{>m�[r��j8�*6ۓ�M>z),pteZSgw�z��˵�%O�{� p�R���į4ֶn��d�'�v��������I��dݛBYP���-9t+�K��~X>dV �6� �1������Eڐ��Q�/�/��hia���EuFs�6�ttt\/(��@�5�/~�E�sA�d%�B�^j`pp���6�P�����Az�래a�> l�V��	�um���/�k�>u/_�UK��YL�	���H�m�5^�Q��7��q����K�S�$�ϝ-H��M������N�ǙE�k�7"�u����ȕ뎓����J�
\�9�x�E0s�5���UQV�m���ꕳ�Gm�#(
�-I��A��o��eݬT��a<z��1����%o���p��sh�w ���6t�{FF��G����$��i����w�ES[�5�{�b�:��;E
��V�����-�J��G���y�`�I^,i*� �� 2���3T\��Dy����OX>���eH���A����[J�`="`:s��)��q+��r��,���Q�W���i|P8�0՝;�#l����-.�N�u\���'��ld	4����եߋ�s+h��x�ro"b�}�e���@������Z�Nc"oJ���A�7��_�����0���[���1���_L!/��Y�MGH�	��䛳� ��Q"��vdo�{�h����$u�Q�@.|_x%��W�q�{w�qN�I~�hM�1����O���d2�r����C����A��M���Jb[41~:F�T���R�i$�Td�����=(�`)��{�
��G����\�]T�:@�����r��^����aPY�LͲ�c�އ�����<�}<<t*xQC����#�!���r<:\Rc��;W,*����X?X�x���<�Pc%.�r�]�F�;^�.�Ǒx��b=}77]�U�y���
n������'�Ӱ�wx�R'؟؋�h���vc�f��Q<����	!fn4`c5̑�$��ʳ��id�$Wɖz��^m]�p(w�GX�\\@�1��b��k�7��MuB�hZ��_qcأ����e��>Qm�DiL�������f��L���=UL �N|�4RgV�������`�8���Ʈ�K+��/y_��7޷{�A՚�����e�:'Eg�ϑ)��"��S��>�tYt`x�"0j�!?-�����V����@�HǄ��x�s�S�ٽH�����4�#2��m��:��j$�J��L��L�oݽ�����"�v��� O+�Դ��My�ɦ���|\�v���q��b�x"��FtW���nA<�7�4��^��]�N�ߨ�(�Ҵ�I��������wn�̧6i�i�pu�.��M�V��I`P�08��H��>�(2+|>��=���;��7��n���N��8[��,�:��ੲ�M����2�6W�g�X�j� ܬ�C���Z�b�s�ъ!��g{ko�����";$r�?�f ~��\�6�u*�JSSS�ƞqbr�İŧ �j�<=BT��U�thb��N���ņN�#�����GL
?ˋ����t�W=/�:n���Ȫ B(7����7���a_�W��&�06�c�p,Ҫ�Za���v��oF}���
�Lqw���)�:2�QZ��9:6�_[[{�`L�~1�,�K?�tw��&AymdB�cfd��R�S���pݦgN�?�x7��P�~�Ɓ+d?�ɥf�|ڂU�}1����SY����5���턦�������W��f�F�jFx����!����tL�G��W�*�PavB�Ѿ�{�U�g��d�(���Svf��n*����뽫ч���F�-O�ǆ! KtKt�n��/M�/�~կ\��#�<����y9��n�f�~��M_�P�η��~oL\ϸ�߫?ݪ�f��v������%��	�d#��I�ɛ��1!MV6�>�Iyԙ�8n蔼�VdV��
$^5��G��������n:!jp������+�r���'��I|����RK�O)�2��>[�4ҼE/���)W�/���}���2�L��
¢
x����]O��8�Pm��Ɏ�\�J��P�8R��S��bp��Kx�^�=^S���6���?j2[�D��Y�eˑ����Q%��_�����g�'��y@)1������6
��xT�x��ݱ~�D/�	��KjW�Rzܻ$��J���j���(�yg$c�n;��Bf��'��1���s�ͦe-��T���8׽�S��������H�gc���5��I_S	a�K<���e(���T�"�{�=?8?�k��G�Ee��,�rI
f�lm��Q�d�;��~���+F���ƪ�Z5|]�N+.��2\A��e|K;�K� w�r.���C��<�a?~SHI�W�Sp}$�J/����p.u�,C�fW*Z;i�(�{���p��ȳ�-K�&��� .��)[>==�FH�u�h%"c��$����y����-yړ�-�@[�k���=�oiy��sf������y�-�z�=:~��:㱧\,JN��;�/�WQQ�sz��CЦ���`��3����{����#Ň>L�{�f<y���_q�����3�x)O��[<I@�D}�z_�4��w����;���[H}�U�.�ۼP�}5e��wjX��&�1#+,DG���ڄK�d��2�ζx�1L��%]����������q����z~�a�R�1;���}��ϩh�Df?}n�����Q':�v��R��)"��p.�q1i�	ͩ��b�J���&N���D	�M![�����~���L�t���a\pZ�h������{���D���!x"�+Ap�(�pY�<�e���<y�dd����9�	�l7���=4U�e@h����#��w��DSs���df^qژE;��YY}��r���u_IL���a�g}q�E���#R%������}8�F�g��|�W����4�ЁbU^̜azf��X��苷Dw���OE�ʏPG�����#�'�v���O�����e�v�2w�����G�ҫ�t����Y�Tf�:MY(uq�<jr�tG��$΂�}��he���f�\��v.�+eK��Ǎ��Tu�G�Q�Oyq�fIC�(�L��x�o,���)��x RA�ٷ���RU��$�^�Hr� pD,���}�%�[�(0w�+p��,f��3^pӪm��E��^M����J]���ݏ�w�Z�ͫo���)C�ٵ
0u�����]�4���~>��A><<<Vb��p�Ly˄��|�t8 ��ՑlG�Rin0������)%�uB-(���ב���#���t��Ru�|���+L�1;��h�ӪaCRg����뫴^����wno2�P�V���MI��k���8�q�"�N��u��sb��bp�}4������yv�}L�$�[��'��O5o.��z��R���65RhYӒѮ|���~2"�o�\h�_>P�_���i[���2�p�\��@��b "�MJ�� ��jU��s��P	�(Y�ʏ�M�)��)���]{1����ڹ��J.M;�7o�c_�X�`_'����Pޛ�&�u񥮎*==ݟ��R�hz}�m@Q0EUWW����/P3�s�p\^��Y[�Y��A��Q
2&H��� (T-�)+9ާ�TB�����SQ��j��~33�G�������1�,����;l��ᛓ�ׇB�~�Ҩ�͗�+�WP��y/��v����Y#�5�.���Ol��Ll�ҡ;B�,2G��܆C�%�0��f���6������S�	/�;CY89Sm���>+�T���'q]R'r�R�$�o�}��[",�s��� }�����U��;���w^�E,p��HuHF�ܲ��+ϸ赁�F�ߢ����<pJ���m�83)��l�9C�]��Y�L�@[I`R�w�uk'��pe��z�E�ϭ��Qb�~+[z_9�癭�?������>���"!�"H��J���-!�ҍHwKH�t��đ.��Н����{���ُ�zԳb�9�kͽ��ח�!����V����&��}�v8T��Rr[/ϴ��f �������]>k�mAro�@Y��IO�f|�L��x�c����s��\��č����Ɲޙ������
��L�oW�{'���2an��ܝ^��XQ����@��ի�I�0=�$hu|qe��
GFN����>��Ņ;;;[�T�=>s�H���7w���P93yId�AB.��9&�_G(�3P�!!X�dX_�*��|s8T���W�N6$<��L��������4�@��N�=NW~�𹽿�Ә��X{#���'�����͟d%��~��	[���R)2/�P֎�Uib��ob
9z�Aٹ���\k���;9���8���׍Π�����n�`���&=���O!��v.�U^ẫm�!v�w�Ls�q��,l����FM�1�w ���@Q2yab5�oo�iݔMRI�r�}�3��'�f%�U�'&N���u- C���3���<�XJ�ڵr��;1����굧�Ѕ�>t}�������퇯#K��P��@�F��Kh�dߥ0���fs��Oɥ#�5*�f%�L�Ϙ&�|�����y��_�F�#��݀������e._H4�Qt���
~~�N�v���?��#��%�w���g�%$)u��3%.Җ���@�>�2�@��ǀdIBBB)e�{��~��e�-�-%-�ee�J�&�%5ޒQ�&R�>0�����ru��_\^�Dw8���h́��>��\�z��U�"�oL�ޘ(����s��&"m�F�v�/LZa/輏"L��ƆzB���11�
�O�ϥޢ�ƚ8y��H�|u�r8d�Z{F�������ؼg���'�S�[�J���m�ɷi:�<z����wJ�@̱���$�v�����u0g�wg�(���d�Eȋ�(CF|�<��Ȝ#pK�.�?�[������(뭟��Ò�b;��I��8�4��YC`� �F��� y�椻or<�LyĶ������X�H<A9�B,	�b��of��߽ٮ����{�E�d�[���վ�����s�׷{�>� E�Nm5ʞ�b����X�`��U=2��J��o�gd_~��}T�k�B�y	�H��R��Q/jy�Szv�G�_�P��"l��cض���/�{#@�e�E
� �{�>M��[��v�`<# 䖺����[l�@s����he}����P�f�7QCwߟr=8މ�{�p�S���;����+�Y�o���F8"������F}w��3��(�I����H��S���MR�-�,Y�P�h<}�ڮ3����8��}>�s��xG���Pkzz쌡Ȉ�����|�t���������n�CE_D|�ˠ��0�HE�u����$�>z2RJ4��bX���jd[����ǝ{�=wC'�����JlP���AZ}W�����E�i�ǔ�B��ժ��� 5�J�6i̓�b�,w�W��.k�><�U�pj���7�B<R�ጿ) DMMMw�����Hd@ɗ�`[�P�[|bo���g��F�?� ��`�������FZPwD�}��m�pm��WzǄ����DPP�߻w-�����1���>�
���Ύ�q�5x��֣��D����"ы�i������p'��s�a��#��,~�P���f������)�%H�5)���ޮ�ܨ˜\UE�H��>j�޺��>>M7���rX/j�d��e��7�x=.�V߆��J�7O�A"�޶����tqqQj'�4�� <�2)����Ν;l���,�&��x��tyKC��0������]�?\�8̌��r>F4�Ӭ-�H�Y>Ackkk���5x$�j`]�X�M{b0|""Q��`@)����00R�����ݿu�Z�/T�b�aaZ��W�y������Y�=W�[0�v�lSz�_�ZL�].F���1j��0H'��::���T�����d��������Z%/�?�\���e�৑�U��U���9���B�f9��}K��?Q���c>��z�����p����7��@�Q*۸��(��������B����A-=}}�@s�@�P]=��X��oy���9S:�1�ߢ�ˀ�l1���Xd����x " �/}: 聓����B|G''�хg�dd��Id>c��]�����j�L����k��.�iK܄Y�Ӡ�ِQ)��o�����m!w��wD��rpPj��f��P$�3R߽	xRz��H1k4�ߠ.�h>!�'��P�e���:�]��M��5�;�o������.�A)�^	C�6�����<ߔ��W�iyG��=�=S4�3เ�n�ˑ��G�0���XqG�VF��R6,��G�.��X��0;����Բ���i���f��7`�u�M˜������[��)�g��xcĴ��`�A�o{j++	&��7�}i7y���(�q��$N�!�RPP�n��D]D �ϽD���"51����C�bbbr����f;�ԯ���*V��.�	�����X��������r25��;hfL���v1����i,����Y9��8�O���0Hw��_�� ''װ��8�������f���"`����t*%wy�z�6֪�g
[H�66,�yn�0��a�^�i�FA��|tt4�i/b��>��|��w
��jA��,��>����)����1!ǃ؋�����|�*(���}�ؼ~�ĕ�K�ϳM��^�Ǒ��0qOL�O�w'���&����w?� D�T���%9��-�F��G >����߃��0_�b���� �gb�c��.�7H�1`500x-.�����+k�xu��U����{����ρ5���'����Q
?�咈�J�NG�ﱿ@�~Y��@WqYb*=a"~sũ�Yy��w�:� ���&�8@������c�7c9�T �ѽ�{(*'��<�Rw�g!'����uy�(���ej��^l�������5gG+��$����^B	��s��)����\-��e,�������Q��uH�����@�c:��`aQ�!�|<���>���e�s��)�T��Jnl���h���񝬬����yZ�9 !�YY�>p����������@��@�zUK�p_^^�ַ4eUiф�j���/>L�����7��c~�yI͢���?0%� _�8j��z������`���;H�\���DX=b�X	;>���<���; �f~�&ce8?�Z|�Xcy�e������>y�Qq0�o9b������l�d����V��QdH21�`Ee + �h@�� ��IZw_8:u��<_R�4a��M��Ұ��m2R����uQgA�z�&�ņc- n����W��Џ��U��{r�e��S�c�!��X=�k�Oo����|ҶQ��/��*u����ycu��(j.����B�����AxC���1y	Ւ���M>����_G���i&0<�����C#���Nŗ3�=^e�Tj���tݍ���b���$2������x��
�<��
2-�*���lox��z�(5'5D�V(��V��֗��EG�W1����m��Дs&H�Y6��)]��G)��g�?�J�'������6v�!h$�̼</06�u��	v�H�\݆���"CM�|�Y}�.C͟*�k�2M�Z(4��4/0PO�W���
ƎQ?6��<`PdT��A�4�>U/�����:,���v��1��7s�=���~(&��활*,,��#��M��_.%T��R���Cו�"wk���p�~�@s
�l�H��� �W��m3eu�.���)!�F�N�ޱʑO�=Z�4�[R>�X�_��5��tDZ9��,����ga;�� ӗ�}�9;'N�K4?����OǇ& ��1BĞ�t��xzz������r�h�.T,$:113��u�~+	~a]�+�6\W�τ��?���.��~@ $���ڍ�Sd��J�,Y&r�Rڰn���ŵ`#�'%����������(5	�J�^�F�Je&k��cn��ǈry!ɫWB��ˆ^�%qv/�{��A�&d���Q0�8��= t��Nw��(�mm��)X�;FE�YyjY�K�/�)K ,%�I�>(ۇ�Q��de=��U�S8Y�?�U�S�:^�?������W-p����z���>c��Qxz0�.w��^�4vU&����H��	�����{=`&��ʣ""�KKq�ѕc�y4j���	�(1�Hf��vO7�~��َ9��*UZ�=�}p��`ra���������]�i�_1F��i �-m�I�</YY?766�"#9e���7,Y��<���P��38��(&�����P���M��M���6�k��s��}@������%�eC��αo��Y1g�������:�
:��
�n�F�j,Q������ E���$Q2��azs_J^��B)o0w��b��}W"�����Ì��*Ԏ����W�z��	
��h�#-�9.�>��م���l�q
m*c�+y` �a�<����V$| �`}��MF.3��`(�7`�n�bs����.Ƕ���� ��Om)���z��Y�K�&���4�O.��txr��eP�t�1@�6f�')!��(� p!��B�Pʷ��)|?FLq�^�������bl�a�U�6ݟzQ���xӉNk�St�/A�	?ොq�g�?�5������k���G���5 h�a(�izF>�>g���>8��?0P8&!�  !!a�ؘsC���_�D�����Ȱ\�R`���	����-���U�V�(j
��|c1��9��m��{a<85g�ݷ���OL�+_���N�[7 ى~eN��C1���н�?`p����G���p��M�H=�¦U͛��E��~��C���� �e������5K�X>�U��C:�G� / 5b�ajJk�U��2EEE}��b�͢�=��ꠊ�J P@ ���qC��!��Q����b���n��p(s��bN��멙l�WD�(=rt��Y�^��V�]��s��w=�/��� 芑�?����IW�h�_��	&��}���{�S`����Ot�⺇.�tѻ,�w^V��EY��<�;F�L ����#���;�;��֏C�t�sz.��YY-�8{Р5��nw���k�Aƥ*5۝���sQ7`����7��K�o�Q\A�2�
�~���{��-1B���F|Y���S;��~�C�_?J�yt�Hq
j�S<5س�&��_����{���Ǌ�O����ȅ�JJ�g>�����Jr�
��V�Y�S �AG�y�ݽ	�w�N��'T��f��cu��$��Ey�+/,� ����OK����(Pݕ�+o��d9�DTD���uS>����I{�Iz"��H�&�TҒY(���d8�*�\�"yjNz��-"\�sk�9��E8:�O��E�`�s|���ԅ	V�NY����,�m��?cK�`�QX�ڒUu-�Iܿ(w
`���}3�g6�^��}��U�	��h�^L{1�xף%�7^�yV~\�iD~���6$|�fT�����J���}�[�y�5�� ��O�f�-�%a�wv%T�Bf�_U�I�j���Ė���a�����
A���~XU7k7����ZW���� @W�#�x� ^�S�`	�z�>))�(Hk����ӧ�� ����L�핿/TB!���0��H�L4d6��	��i �V5��<�Zq@�%G3����xϰ�r��9x\f6��ȕ��W�ߣ4n-aU�r��+�}��q3ff�o��n���j7�����4f;j
&՝������o�O��UU~���A�E��c��˿�/+9�i��'�#����ӗ. ȗF��O�+)��_�V(���=��-/O��E�y����UT�Ć#Z�?���~`#� ����(x5�F3?�xBvp��@� 8�x�xV�� �#*@0!���d
Y�P���*�<�SU��4�̗�D�hR�U��W���v������g,��;�K�#Z�d��s�Y���^:r�{O���^�/Ŭ��9U�HX=y-�}�q�Ipt��m��u��rJ�K�xq©B�ʐ�/�:�r[��f,;���TtYvJ���	D���f�ܮ#���΢���-s��F��no�b��b�y�ʺ8y�����g5�b����jdb޵Ї-ɕ,��=��ő�4�e���Ԝc����/\�NM�׎�~�Xw���?N�Ǌ��e����@j�t�Ç9��"�A-i��Ɔ�D�#C��:��ĖٞHz��u�����ݜ��b$��F^?#|Ѩ��Ja%����)��#���uU*�YŹ�<� ��@Ǖ]Y^�	jyG��iϤ#�[��=�kB�gaGs�z�2������������ǯC����pͳ"����˓ob���k�p�� ���')�_��������\8c�Zh��p�;i�@.� �����V��`�&�k��1�8hw��ƥg���n�ӆ�1�n�;�y�϶:���� ̭J�c��_C��@pyκ�_k�U�(bp�t|r��F��f�6///5p��9�׭���X�뵷��I�ۉ����W�Wh|�b9n6?���p̪;E�����}�/{��UޢK�L&��&r/�I��B�tw1�r�Z�u��>��T�ecc�@�_��˪�R��c67/p�
K�,+��U��(�⡅�|� <=�<�u�I����S�_�M���D�"W5]^�
k��Q0���i4������>�劙my��9+�r���	�:N{=,�'�4m�$�{Z2�Y<&}���X�������cƋ��ݳ�n����0?�|<y^ɨ� ���mbbB�E<�G�X�+�=>��6:x/mAMʐ��i?y)?Y2�I=r�I.e�B���lIN��Ą 0�ʥ��/�^@�߾���-�pn����t
��;E�_W9��@4��71�IK'/�ep�?h���cq.JS�9������.*Þ�#�d���V\���6d.���si��ۆa�R����c���jf����-��"��#PPQID�ie�A�S�lU��W�D}�����i<���kg�/ق��(��/�*�=s��ڮ�������B�"s���z�M��/:��ggS���m	Z��=]�|5����J�Er��2���>�u�S���ٍ¹H�����7+�\Ը-�B����j����˖rr���a�,.vK����� ��=?���, �z)+#qF��-6�2� ��8��-��>W^e]�=��h�b��w]�,�w�-}�8V�q������v+*
���>I�<��X+��������d_X��L��6�hf
G9�����ŉH2>W�E�w�\�sC���
وI-�� b�+ ���"x*+��9jftMT�Va���4>���tc�g�kW�V>��
��ֲF���C�(d<�a:jd` ńOl)fk[���)����D�=�/^(���vq�ǃ�x�+���}A^���ҥ�ei
;E��"�|K*�)��˻^�����R�zjQ�baa����,���o�܅i�����]\N��41�}�&0���Zɯ&n�t�^8��Ө������u�!H��cV��5["�ey�����о��?>�}e����w��T�/��'�C��-�rG���O�Zf�ΎVl �c�<:^$�w�X%7�l���y�k`�R���]O��1RZ5�J.�(QaRTTF{�H̳�����څ���^�ac���ngʑ�A�P%zib���qP���ά�Ĥ�~�%��R�N��?0���=�>ZLeF��@$IaR\\ �2f����	�Ň��AC�M�P�5�k��ui�iFԵ�����.����٧1JfI�Ne��3�*��J��s���~��ھ��VDY������O�H����Y9`����u%_���UTLg�{>#*��"�o\^L�t:1)�`$ @
���:9qI�� ��1����H�Pk�aSJ|U276�[)��_]5��헥������e(���ة����x���E+]@W����VT��0��E�3 Q7 ����1(n�o��QVj��/G�=@�&���}�/l�����6�Om�T[�țZ�W,� |
D/��7�J�k6��X�_� Hs�{�YF�%�o�����W�f��)8����r�^�� a�T��4ŕ�
¡�6�G���
W�Uۀ�D"�x�9+�,��)|�nUc���?,���4X�eU��䝜�
4�8�k����|����#xv����%0b_��І��y�j"����4
�L���RVV�xv���ӷ�$7�i{���
�N؈w�4Љ^�E_F�����e���m�Ћ6Z��7�F
rs�=1y��Փ��!�`A�����r��hFr_���nU퓘���{^�Vwl�0֔���426&�@��)y�3퇚2��vL>\��d��bBbs:,*Pƽ��������V���7�ǖ�B���E3������R=ǥ��_�ж~����!��m�Z�Ҳ2#--�_g������ �:3
�
�N�Ow5�Kњ�YY}��GfUK�\�G'�q������݌5Q�%?Yj�NC�@���*�񔍌����"�e�,��T��2�8D�K���w�ხv��㸼�f���=@d������:f��G���d�%X�22qwNA�v^A�$dwCì��u4I�K���[o��hH�ք���§`�\(���t�A�ոu�(B�)���XN���4���`b���Cȏ���G��H8mŠ���S�ת���N%Sh�ԯ���~�ӣ�޼��ap�I=�&sA�"���ĵ�CG�,��u�z2��)<�PV�]��IWU0�n�tS=�1���&m�.�E���U��������
��D3��t��HS
]��"�M���2=t�2�a�_���/����f�ꉳK�7[ld���;�ϖ��V_���5iv��Ә��x\��]NW4�c�$J�G4�^N��nl9�
@n�� �oĹ�5u�3�e:�U���=��k��w�B�2[���UnT��UpL�[���6��,�H署o檽��3N�ܠv��$���b�
��"т�9E�Gi�f�:��x��,$+�F�mk�Ҿ��WB=%�s����(x����[Ps������F�.3W���u������A͛i`�-S��4v���ȯ�V�ꡕh�"ٵ��F59�����]Xz�=W���VT�z�qxT�$�> ���^��7�v�\�bgU/��I�p?=�"��ʛ_r��n>8�$`�l����ez��O����?�&AH�7���0��vg��k(�j((G�U
H��+>bA �VP �9�}����f������u#I<�	��g@gdt�gH�ONO�;i"�M�B44�E�*��q�[YXH����f �<?*8_���0~���-@>
g�)R=��:���}(���	 -k��'b(W�P��WӨ3�ݘ��*bO�O�]�J���U3~�@åm>�����i)��.x$}մ79�x,��b�|G\m~���=D��y��UW ��1�����3̑���(���S�L�����
�R��QK�p���G%.:�5��	������B[��̤*�w���[��u<?��1�Vc��1��';�K�4B��YLYÑ��7���p�Fr,�]�	���[+��*0��ԫ��頼BH�z�쨪+pS�)���O��Jz�s!̓}He@�TTUA��޷��b�8/��w���p�MN )7��(���b��xu���zg�:��[�]��b;��E�#����遡�����m:Z���xǌ;Wj�T�s�g_�"!Y�����	�p[�Nގ��e�<�Z���kk���\ ��њ,�H`i��E;+��*...MƍZ��sl2n�'��~}?[G�;�G�Ri�?ފ;�*0s���������<%��,W��4�Y�Z�-x<�ŵl� �UmwrF����2ט�{���y�20PH3YJ��d��)9��7�B""�>�W�,à�>�?-4�+��d���W�>��x�.��u�W�Ѳɮ`��fc��4j�����%�4�;����N���(��Fff
\��&h�&����*@~�T���h'�%����o�bl�2dݩB�y?���͚Jd������&�8��s���^eR��j~��Ū�*V�Ek4��2��٣�`����,PV1. (��k���R�����Fp��ڿ.3�$Au�]�iK�<���w�<,A��U���Q��"����_�����5@R�p�3A��z�a.B�x�ݹ:'G�x}�a��mzͺ�F�ko����Q���M?��@�%����N���d a�j'�pIL�w��B�H=a�X5i�'}��`L��w�h����5�t=6�z��{��B��+1aS��
2������ō�n�~���|ౖ��F�A��]��{1)�}�+y��55jyyy h�V@���{�����WPw��a�Ǻ�g�������v�,�	8�
I�ɊYh�v�{��~�8�\�
��$�PS�Q����{�@��W�޾y�������5"2�2���xu�����(p[�� *u>�|ՖHiT#ΙcC�FE8H�a�����d2fj)N��ܸ���V�;S����%%_��X�A���:�]S��@3ն�����0�ɓ����C�5Pj���ސ���w�sܣ֥���-�_]7M^��z�3�R���ۙ3�-��]�ܪ�A-��L6���מl���+� W��ӫ:��#��><�@�"�����w�eM�fLh��5�� 4�/	5�]����$�W���d!_889}����奤�@ǣE�=;^ǜĸ�9Rj�_��:�?�9	ss�h;�Zb��]�}[����G���������i�{C*P�����2�MK0-���Gg���ʦG�}Y	�0���[�j��ϔw�T��0i�S]̤��(� ����m��b�5?/`�M��98�'�-��3w4��G��, s�mK;;�<Woӕ	��7y"��Gם.G����ʒu��PZ�%�(�7�fD:ChK�0�����������Q�nګ!����߿���Y2���剛ן�m &&4Hح�E����#�*d�qQ��f�Sv�@2f���RN���A:��Z��˩xy5��.�M��XQ\6��P��Oh���{�����q��+�s���v�v�J�͠{���q�"��J0� $����9::����i��fP���D���dZ���Z���z��#�ZE���U��+d{���b-�r�0�C�1����r�>K�{�P/Z��Z��� �N�L[
���+��ؙ��j܄�1bz}yy�W�nw"�:o���o�#_�*a�<mM,v��@*�@���[�gK�K��T�`7�Rj!ϖ̯���Ԓ��e�����ި���L3=}�a�#�t��Q�Rg����5�U{����MH-�ġ�okEn���&X�%�e!�������ْ�ВF�2�Qt�Q�	�"D��)��hB^�t�3ri>�G0�dXx���>/E��[��/���!�#bI����**�+��\�D5e��d����،��b��I�Y��2�kU+`-�rO��W:9����k3���Y_�u�zWY�XW�SD��;�{�x2%����V^q�r�7��#�(pqp2�r�q���J��,���-@����AsQ��-�fލݽ�,���os=�"��H�ϰoEv����xS:�ϴu���N��Z�#�s�	]��OQڀ���"Q�-�c�I�ÓӺ0w����o@
-$:�/����g@�����]��?�����T�}[�[b���ʶXy���F`Y1K*f2O�E?{���?%�g�BXׂ���%���h������v��q�r�>�TC�W����z���Ԁ���JM�:0s�d��f�n`�s�ׄT�d�LLֆQ��1,��h0���ɕ��N�����8�� ��7Z8��͑IC�n4d�����ȗd	:�|�C7�,q�g�Tp8e����"  @CC���]�g�.cl�H�$��p1�<�m�Ɋo��W��Y;���P&m�[��><���.��:#E�U#^��H�k��-�'� ��b��VO�Ji�Ւ/-��r��l�:l8���f��iV�o!*þL{\\���-(�.����a����Q��ꥆ��%�=L74� ��q$��
~�t�y��蹜蟂�1�9�����T�SU?�W4k��%"4?�4O�.0�+3��c����~���i��&�l��i�P^.~G���!��~0��Dfo�7�'WUqd�^%�׿7�E���
���A�g��֣*A�%����h:��^�Z��0J�uI�!j̬<\�Ack�U˚�et��z蓌1b�EP S<��z(��X:���r"h��ړG���r�����j�V�wxH���[���xw�v���D����V| R<�`K�4��^^\�� \5i'��-�׽��3��vE��t�d���dε
>I���+<N���k�Y4����VH�E�O�c�!����Zr�{��RM��h]vvv��"���D��+(D�h�}t��ԣ��� ��hn�����Փ\]���sJCMF{R�KWƣ�vFp/8>T{\ٻ�<h˜o���%P��:z͚x�%�r��=�v�N����H6?�a ����4e~:T�? [}j��pّb�����}�O����e�*���n��7��?y{��hX���i[�YmYʕ�*�2-�''!x�z����vo�֞�sqY�$I�$�?���YZL�RTi��׏��~̤�qB�����n�����$Y���uԋ�m�F㎖��{�*��ü�	L��*�?+� 77w�w"],����,@�g:^M��R�������|0W�F��t���Y��*�%#��#."St�ۃ������:S��K���\8�����5�������k��67<g��pm:�rǓ��Z8::��o�X�h �h��T��T���ռP���c�ex�}_������H�����wnh]]��� -���P%DOO_d�*��BD��X�� P`>�|��� �=��B���wFaZ��n����_�Z#S��J�_��ț��5������{���خ��f�^^^4tt��=iO���3:���D	�j

�fgiU�zu�4j��2* �8~t��"A��L��Zہ�����~�l��K\�V( ��i�b�}��c���`Fȅ��R��q��G��v�f��og�/B�Y�Ӿ�w���\e��F���`V���Ȓ����s�[\J�im��b�(���礥�SPP���������@7� ui:J��/egW��f]ee�ȏ3f�`��n�������Y[Q�ӝ"-� Vm���`r��<�˥u�PhvN�M�퇙YY��l:��bҗ,�a�?�DU��L�ǟ	�T~� �5O�T��n� �)��:�w=��٭`����֥�-b�l�|�}��)quyaa_++���U,h|�o_�v ��&��40<|���/��)sh�z�����E�?M���Cj7G�Q��ja[��ܙ�^ǏH����ŝ�p{��tS�hqq����?0ǝ�@���e#a��%6�|u1˫$�n���k+B������DO���q}��x�uK�4��6"�ێ�Pו�c�>~�<>� �?ߙ ���ܿ�	�ד��5kS�J���rҢ�������Y�^���;�E�2�'���֭����Q�q5���/�v�`wy��ĄX#���/���2�����2�V)Ě���/����¤�:_��#^�7Ş�6+����:�g���ǆ5_��z��"HX�i�|O�����n\�_Y�}��g�f^�-��B1�7���v�%��H7��|r�yLY����&_7��l��}v�*,���#K{�WZZjğJ�s% e��ֳ�d��w�7�����7��YlO�e��X"��E�䭭.�eg����	X>��n�Ꞅ�ǧ���~�ғ922��ݞ�g~��ʐz�?��Y�#CI�X��1��������p��&���׀>{_m"Q����^�-(f��	L+�v�7�J�}!ȼFFF���+��]����	������4?WII��y�3�rw�Y�ةli��LDO/鼿e��""��z��ٞ���r���� FB�$��n{6>�=t�r��ü����L�8ρ���Cۋ�	g-
m�r�Ȃ��$ ݄C�.�{q~��@�4:�a�DbX�,������C�	���IÅ:>f5��>�פ���a{�^t��r$�	�7�o��E��	�.˯�����p9��>��,X���$|W!_-�hT��oSi-���˿s
���3�烼F�+�b�˫�j!�>�-�HY�WU&?~�|��Z.�Kc�,��>��pXH��������24�F��X�RI�sI<�U��Ŝ��B}�:�����\{��j1p�W��4(���&����uj��͔�� 5����Y�E�&�4{:�pҹ^�Eȥ�)(�OY�_��Ž45�����o�r��B�v��a������!�u��1[M���:����?�q�=�Ӭ���uc)�##"��!�� ��A2'� �~��rJJ���xtJ�ޙ���0O�=j��%���f%)x'!�u�U礁R��j��Gm�(�(f��5�4+a9�o!�CM�B�����{�G�(��k�����9 R%M޿O��w1����[[[%�K2��Ur��nt@@V�D-{���ή�r�q7S�� �[F��ƻ�1j�Fook���LJK�l��Y8(^�-�������d��fN�ن��YT����"vA���q�n��v�/��q���cP��\HI!s9,#*�QMmX9�յ�L-�6Z�{���,����'@��տ���)GR41�)(�[��ܑ&�ֹA8 �I����`����e3e]���R��v'*Ǥ��$����R�
m�;���```@�P����/���%��t�õ�J�B������C�
mN�R?��q(��G�pyih�8P�_ժ��S.d���8-y	va=jC�cBӄ�S e�����S�А7�;p��&" ۃ����w�p:W����3���I���8�c��hH�������Ud��w4�o
��v������yA^�}�Uo��>8:9A���/��	c[�ݟ�%	�j%��z@^qs��*���Bӑ�_"6u��� �j���V	��p�J�`�E x�c����������5?\Ǎ����3L�Ra˟��m���\B�מ��� bW)�����"��$j�9��C�����Ы�������tUʳ���F�
���TJ�?sV���TJ�Q�%�`�U����� �wJ9ͺ��4��
d��L �p,=�V�'�$P�p��"�@��HK�u��܃��0>�O$��bqz��W-j��)����{��t�t�_��YG9�՝�����/r�I98T�/M5z��(7U-T�1�>(6!ДDp���Ǫ˷���Eڵ�3�P�A��c��?݆���iYHH_zS7.�rK����c+F'%o����\{����vM*��m'�6�+3?~�Ḵ��|�.�G�1���-7x As���l�^��]Q����;h�-�Ɖk= ��`�L�o�--�UK���Pr�fWw=����5�gU�=�4��#��f��p��r����Q6jI�����!݊~颢�ۇ�	OH�S�h_���N�r�I@j0R��?ȧ�w��/I�x6ٮ����-��g�ߦ�@��1I6��*���,oo:�ܺyq4)�Ҹ�� �:@��L]�z�X{0�/�r�bL ]��'~�� ��5fS�[B�x��t��`KZ�l�el����I4�S���(Y���[���*BB-��B�B�	U�9h��������7���8�I~d���15Ed��jh$�Vl���Ffȏk�yE��[��3��(7�tx��Δ��	1$gv�ڻ��� a645�wq����-�[�P�l�u\���y)��؛�p�ފ�n�d���0(�v��	*��X/ I�j`8 ���Ը�yÀ�𸱻��UP 	�Uf����o�R">��Йgna!'3SH@@`˞#�ĺ/]<lr}h�ɧ�n��F��8��qzW͢������^E�6Ə������bl����M����Ms�7`Y���/��!hg�S*|[m�nˁ!���D�[ng�DF*��+-i��e���y�p�e�8��k=���5K����P����(6����Ձ[�@��2�$��O` �0්���~���4,XT�m:����@�cc\Fn��
�I�g���MC}��5�飴�:���;48�����ᷫ����{0�{$�B������	�xIl-~��Ƃ��	<���hg5����j�U�M�I��瀯mE�綷�w�����A�U��v��9Z���]^]�377��~|_
<�� ��̟�x;��w2T����SV�Цk��H�:�o���y��-ؑg���ْF�ϓ�����=�Z��jU�E���qza@�C�sP�bh��<�9G!/������|�ɒI��>��R|a�/�ƿeI��$���(y?V�� �ѝ���3���P	��#III���sVByQQ(l?.H�x���4���8B~@�x&���'�Y��<��)g6�bJ���3����]�����l���޽���-""x��v}"π�&
���i� 1R*���#5�x5�?t��b�p��<��MIh�t���n&%���Nh�kpp���k /XY 5䰘r��eβO��xps��l.{�^M��l�* a��� ����؆�`*	�6���]�����»)��I��hwe���0��a�N] ��`*�Enx~v�Rn��tq�kZܧO7q���Y}��9�B�- %����
'��"hց����kPA׬�9 ���{��GG%n箦�u�@�Ά���-���g@��K/gl�Cgl%FaW=�Re�\���q��[��)�|�Ғ7�Mn?Lk6[W]ҫb�iW��; �H$n����7����&=׹#������)���AR�J�RQ�d`UO��r��$�|v�V�o�l4a7܇YoL�i��첮��e�������t� (R������<����h�	���}��%�����N$B��'�ru��L~�q�~�W����^M�g-�H���p�32:
0����X��l;Ɏ��6��V�䝡��\����0�a���y���
*%�����J��I:�
듅 �T��`�ѳ~'Gǝi�GP��g=$�iDq��d>�����I@�w%��Ot��H�8r��<�ċ_e���p�g��̨�u��on�y�L�=mA{]���8�bG|e0o��b�[B�,_�O 1��6��i	uA==��溔):k� �AG_��w��v�e���fgcc�Й0R�Vӣ��#:8��Uez{ߡxЉW�á2�V�w��%ҢU���|ȡ`))z>]�p��G�g}��nb$�{��3�.,X�6:xN��$f�i�xe���]�n,����͖G��P�l��zuQ�:25�R��)�����Eg�����`����������X���ǽ4�^1�1d�z�L��,������+��f�#�0�2S`{jZZ����(�-���3�r<��_��"r�邱n�S�5E9�Őw��K�"I@.J� ��bj+Sp/��:04Tъ��ϰ�72*D���2kW�'�ګ4�zy���V/��ٹ�^ׯ� 409�軄���mO��E=G,.vC�j41K\�2b��+������>���T���P}���%Q,Y
b�R��Ԕ�����cPSȶdX��c�o�Ru3�b?άB��'UIߥ��p�w�˶F�}!�2^>\�Eh����Y9�<	 _������ͣc��BN/>��سW17�����srrv��pȘ�+���)&<z���c��6n����
�����QXA`@A`W	i�	EB�;T�:TXBPR�s�!D��a:��� ~�g�����}�=�\+��k�G@�Y���u��Nn9�]s�yGA�2�vonA���|��rF(���}�!��'l�rm�B&��+f�2 E�{q��&��ۋ~Mj�o˺?WX�@7��q3��V�� ����������Vj���@��
b�c��+<@-�m�Ėp�N4H�y*T�.d|6���
V:���nn+_H�\��q���\*;�E�C��w���?5c*���� ��ǧM+|@@ �/y-���M�Ha��"�;��	;�v��o� bf3�!�/�v
�liyB+�k�cU � %�4��q�S������5$$$;�#���k����?䈖|	��q��y���Þ T�7�	���r[��$lb�S6��5�.y�t��1���D �M����9tV��osW�w�.w.{=�(٢�_��@k�[�B���q*��x|tJMC���Bm���ZF�V��#�k	2�3����XĹ/He�t�(9C~Z��i>����� ���x����� �iB�e��$�����\�q���+��sN���{?�%+��)�_b�ٸkW���j:/�+(��!K�ń>�=��%6��0���a��&��~��Ϝڿ�� � ��۫����'��?� 1Z�*���I
?�؏��(ԭ�.�p	~~��z8���S�:�Uq]���^���G��+�S��ώ��&�WhY��=~��rs)�����u��hu�+�s-`'�.h"�%��W�T
��E�F�N��OGЉB��I��$e��П�$��dU��ma�%���@��͸�{M2��CPm�[M��){g�h�i��W��Q��@�:.qtT��TL���=vJ�_)�k.w/#d�s��Ma?	b�Y�dr`|�-��%q@�@9��kf�h����o�=�g:\�Z����Q����]ETW=ڔ����㺘%%��珃]o���|�<+/�����eQz��㛞~�ƃH�˵��<�Q	�ѷ�Ԟ9�-�U�='&��9� |�@՟ W����p�E�=�vhv�Tj,�ݏ�'dA���A_�S�c��Rt���g�UH�I��e�fݔ�h4�ȿ��@"
�B�+1��_�I],Fh�bq����
������zßI�HC�!��.ۋ�c��\��YH�ɵ�R� �#n������[���&C;�����mAپ#1��ֲ�k@fj+ЍѤ\�c3�V  Y�5��;���;� %�\~e�U�[�x��Y	(�����}y{�ѫ���n�[��9� R�l��FF�ம�a%F�z��3���sF�<׫,���
�(����+-��/Ҏ�|�/Kc_ov;��ڛpӧ��|`��h3E#^�ͤ��\��_��m��azt���.]2���t缴�mj��x^��QHL��(}q�UD��x�ɳe��(�yG�޾��N���_!���$0 nO~��ް.U���� m��/]��q���Ȭ����Xf�X�,�Zl�[		�\����>��S��Ijkkc����N%��������K{�(i�2_��x��ˮ���Ίt��u���|Hq,M�.Ӛ�9������� *xK䤜S�)Ub7V���a3�D�A��X����˨ͫ׷��ѝQ�ݓ���J@6�AOx&˿�#Mf�9!��yu��-��E󮯭�9��(����~	6\�k�'ٗ"� ���fs��V�8�t����l������<ɻ�CVj%SXQQQ3����|'�ml5<t�_��N|��YZO���������-��kЊtY��jeffR���\�J�h�W��̭K_`�\m���Ye�� �0 X���h��B�~�����\�r*�W�QW�܎'I����}��m���'�vdm�f(����J� lY ���j4�k���Bh��\�|>F�K���v�*��W�Dڗ`��5W�{�����ņ�"�����;{{qU�_����W��h��+3E���%tW�Tb1���k��#������_.���A~�����z}��io�y]N�OV2z+V�%�M�,�9�sM���A 
�� 	�~�֠8�6---N��Vkv�X�p	�s�K��U�$��⻯�6�.e N�����"%%-��.����T������\vz�!� h�Qh{��k�ϵ�˲y���� ��jۜ����u�������*�""����Ȏo^,8!��1r����5W��U�6 [Z��������Kz6QB6n+ ��#��ҫ6w(_��G���t5�7X-_��PWW7K�N;Z�&��>�>�\ᙙC�M��p��D�����-��i:�}�����k׮up_+2D�,?����c��D�hlUdd���Oz���*�@��U-�A}�SL�/$�멧�G�&���J9��ը�����mY��|e��쬠�b�< _�F����o�g����7���'�m���҅�O27�j�xԩ��>�U�X 6g��U���t=�-' P��ҫ:��.�~���U�΢,��������..���{��/���N�^�_@ @������<|iܘ�s����0�TĀ3̎��/�|�{-��w�Հ���XŚ��ug��nL0�j�/:���h|7"���ٝ�:θ������T؛.a7|��*�^jD��of"{�h��O����VV� �궯A��?������3Dw��(�R񸸸䥧��8��kP�?�7C=9����~
��: �u���|�-��}�A�e�!�<��0�� ����:Sⵉے�r�ܧ.����rv����{�����sN���[�l�G�tc��c����'��
Pe�jM<�ʣ��R�i��6]�}h�"m��T1
m�d�;�������L����}���tͫ)��.=�~2���) �k���Jn=�/(�K	-���o�Tf5��,�S&��a|~˻�B�7%C�4Í�P.5p��&$�g��UX}||��
�Dv.���C��===�8e�J)�P������f��Ѥ�b�ԍ
�q��_D��əW��m�����ӥ`������,3�'�Xb��9K\�I�����M=�A^����}�<�c��� �C�\zE�����Xj����=|����?K��
C�B�/��3Z����x�V� �%�����h�P5���ik�4+�2@@-��X��;!l�#���#?~���h�?`YF�����L��xN/Z.j�[�W��rF�ŭ�|nx�^R:m�,�U:s��̘�Xx=�����Gx�w�������u���bK=���/�m�T��8NC57����1>ᮁ��eu��\���>���>�ap�tw܁�,Tx|�\�¾}u��P��u444������`D[��;��t��C�;k��Ĭ�i.ĥ��-���@��l����g��Қv�#a�%~P��}%��>�NQ���o�'�O�p}mL�̶ۘ*r������u���PϬ��$��mƞ��� co__AnnЯp~(��{�6ŏ�Z܁�(e�$c��g���;p����b�0��@ 	խ�g]N%����i-[K��ד{ע��Mx��mu1��]���"+�"��O��:�<V��"�R%��yg�EJyUs���yd�t�ߜ��x�ĺ	q���kM�L4��[�STȳ{Z2����Rq�&+Az��������e�~.{��� �t?��ث������]o�
��,�Ғ�D�/@�b�W�ӟ��l��~E�C5[��c,�������F����ކ��������{�m��
x��M��e�k][�Y
L��rG�����w�~�1�X���8���<�~�XSǍQ4-�BlO���N�!H<�f7n2��X>1!�+����C��	�6���������* �%�iR� ���xyy��=(?j|���.�N9��g)��bn��?�A�dr�M|��n$�8� ¡��Zx�[Zק���]����C=�Xm@�L�
�g��t!�J��e�_���y���3I�� #,�
@@-3�����Q�ە9���bb���,�5�i���M28/���Tm�=通����&��<��pjq1��H�J��UXZʝ�����p���~s@3E:w���n\��C�߽3�Ϡ�D�vܾ�C�x���A!�ӆ��Dy��Z���l������l�ΝV��;`9Y{V�D��
�	�FZ��yb�h�{��4�(���M�~�����)@ 䓓��ի�� ��6M����	���O����j�?~|

���
 rc3��S r�B���1%h��{{�r��>���z����F2�w튑��@��$�|�q�������4&�SC�V��l�p<��ؾ��Rf|�Z���9�eu�b���d�~y���P��`�A3ʹч� �M+b ������D��y��U�ۏ���koEў��Be�y1�����=�Z���@���(�GXT�ֻ<_�K���$����S�
��b}����P������)���N�f{�s��
����6�-�V�	�{�`R�X�3���Կ*��s��i�'�r�T�a���W�u��j����s��RTVnn�H׸���s�j?����tܦˤ�'��9Щ3�.iz�ȓ���R��K��W�=���t�;r�A�΀�؜��5yd��w���9e�'�$��,�������r���ӭX'�T6����W�K�~�մ⹁)��m�MFG���"�{	�c��!��/�	����|�_�,lY�u�Pf�+j+E��ת�G؍il2YGCmB&6I��뉩1 ��f�bs�G2�	��Ƭ�E����TU<���^ ��kL[��w�CO�<	hȮ�r����p��@%��5$����Pg&�R�R��Ï�L5pGM�>X\Q�l��cW�k~���9�-Z.{xd�"�|��
L�`� JB�E755�ހ�nUp�s��D�L��I��zL�h�q�~ )���E�?@��	�
�ק�0���/0����Ⱦ��a���\S��Ʉщ��Z_�|�R��^�g+���a���o����mf���q\�Ts����������t|Fcͪ�55��FC���G�Xo��(yJ �1���IɃɳ��~'a���������	��p�M�r�` ��E�T%������,�gE'ם����
�@�p}ڴ����g��-��d:|m�'{	F⟧�jj��vZ���45}D���2y*��G*N��HFF�Y�%�d0҂���ϗ��m�lVE6�I��<���A���#����~LC��ag ?�mG3@̳����7cK����&�J�G!Ղ6�RdVJ�͟��-�7F�,��J���r��ϊ���������\���4��K���Ю>>���;+�V=)��B�bC$�0
�������)`�Y[���T�*b~;�;�ד*����o�#��A jU��˿�h��E`c�y��݃����\���rp(Yu��3�{�4�@� ���o�P߹S7��~?:��v98��"�������;	h��?�ʎ�؛= ɺ���i?���:�S�V�_�����b���\MP�X�ho���	��ӜS�� ����wG0r�sPx��~J�����+i�Ny�C������A�{��6���m�@WAe��So�n]#d�P�Kp�t6zx��>��R���J�y��H,�{Ǟ�d&�9�Q��hM|[�p�ЧBwsZha*�mmm����r���R#.v�sѧ��T�0�� ��ŮM�e��Z���]�J�~NuI��������&'��O�]#�b���eu�GZ���K/� ���f.��چ1�V�t��%�����#�q���>.����#i�V� R�K�~zP�t�Bsj���Qs�ՙ�D����gb�zz+-	q t8��<c������%당����_�jr7�O��
�ܘ��m6�t���0�"�� �g4�!DeƉo���u�������%��m�;�iil�>^`ޚ_��C�0IZ�u!��ֶ��6�뾚�.��U�k�BJq�	�,	�����>jض�F� �Mջ,�SMZ��K"ƃ?��U�"Ϊ���f=�Feo�]� o�T,ܱ����8�|�|�s�s �l�nE�;���=��-㍫P�����4}���V����!�N�ZG�CϪ�)��q�A=tWo����0)5F�j��^�k�/�N��A��6|y?�}��.���]3g+��I!��G� ���d߄��& 2�d�/���}���3<5�Nq�=Q%Xw7�8�ٛ�w�և���O��6�
��04���oBB��	hiE:��_Q��ʑ�W�Dj&=�W�%���q�2���ߡD�9G!9�2B7�D1#EW(���~�� #2T�o�	܅�
���M9��!򖆏���I@^�S�ݏJ�Ee��M2��7DT��A3���հ���P�/q �`�����to�\7���:r�aKDUom-�tM��rk�̖��:L%����
 ���'��'rF��/���u��Gwɤ�]7l���zyii��A:& �ol|\^ ���}[������/��PNz�'�<@	�p��/���]�:C	p �c��GCn6����~�v���xI//��|e9`��A�P�j�q�Q�R� �����%6�s��gz���\>�txP>'��	D�4yy���cW`*���ꛞ�w.�oI��TP�=���h��Z�D�tYHA �J���*_��Y����#j��'M�->c����m���V�����G��H��Zh5ED
z��м��˽����e�e��ֻ�%�$�2����2W��&3J�CɇP�E2Z�,��TBR��uIWO��S<�������ff���wP+���ܷ��&�����s�,�����2y��w-�x���W� �]�q߆���jƋ�5y#;����o��X�_&$$,����0��o��jV�ag��@��5�[�
��><q�D6"5�$S[ .�ᭂz&�T��o'l3~���$���R.�����XĽ	�T(S�?�j���'��!"��>����~���:9�'��о�u~�*��[������]k0➜��{B���
9J�"ǫ�����Z�����.�w��+j?0�ΰ��o�@P��|VΠ)��p�ky���r��wtxSխWW��]���X���r�mm	@�QA)��Gc�J�#W{���~ǸC��&��'n�8�����U�8����-�"r-�{��׾��&��៖�gҬ���r�nvY�����';h�=�GYZ��Ą5�D��$ "	Ll�J�����E�
b\^�:�n:������Q��笢���=��N�i��33��z�>�ی,����,)w���2Be���;�_���@�^s]���dӿ��W�t	or�%��C=�(���q[��蟩p�o�C�lBb���Xf�%(*(@�����m)	h2� Iy������l+�"�گj.O���ꏡ��S��/<�S^ {�l�U�p��i9�^;a�#����I�����*���F	 -��1���;y�c�Q- zɧU2|�5�1����� X�&%%]��G�-{������m4]!����R2<�_���dQ/-�$	����+ ����:89�ػ��� ���ɛUu��h���2ޛ)x�7��4v�C��������!�?ۡ��3��v+���\wu@��N7"V�|��Q(�u\OR�t�IB��Yf��0�"��?��$P `�Ag�7Jo����I(���B��V/�	%����>R����E�6Q?#n��T)�o����|��1Ҷ(��6���*�sobW	�c�*�^�ܣ�3���e�<'p���aM?����bW^l���#���3�S�7�{M�ԏ��݉~{U�Pϕ�V��n�0G�ޞ��C০�{����:���5�`�K�Fj�>�])�n5��p8��/������%6�* -w֣���,DS�x�+.�G��E�w M�W��e�MJ��Q���.�(�E��w��ם��!�����-�����	hy���l�;n'�_`nN��ןN�6(���GD�<�K("j�_ ����W�;�ƅ���7�|u��u�5W*d�VπTw-1&S�p5�P���ӣ�Z%0�>e֓�?���ho]�+ ���/��AOJJJd� v�8�D�JN+��[Xu����9[U7'�g�.��&܀'�h(��_��|r�б8m'p�T��=s��,=/�M�<>@m,i9e-�l�F��ĥj�`���Z�;�]���dVc�L	��W���H���C�\��˳�#'��s��y=�+zQ�zg��\�/	�f�s!�}8�o���Z�Ǧ��<]�u7S�s_��'���O.���եde̬sv��eX?��/OZ[閨�ϴUWd��8SD����(�Y9W�ڡ�h�����
�8�\s��Qy�����dd^^�pZX�hyOr2m�.n��}�Qv{�Y�X�ʆ	��o���h�r��:����_%hԕ*On:�X��I��^���+B���8�Z߂��ƴ�J΂�u&aq��s�!��z�(���^���4����\:P�R���W>��y�/��6j�ebbR>�f��Ps~�Tj9�~5��(:�N�����ӡ菟b?~�Z޼��D�Ip��bi�N�"$��߼�l�s[h����>������TP���[�b�4]���X̄�ƠG��vla_զ��y߇�'4.E���?���m��.��ژ����*�z�N�(�����c&Q�l��9�:Z��&KT~T��1�u�f��|c���P
�-�������+�=vJ��c,���dTT���	<�cy�W�R^���yj�0^b&¥3դ���\��p�YpEPh�q�6�NQz���*���&�#>11{xV�CQQ�������On��#,L��������"���´���|[r)���������=Wk��s�|�䭭�X��Ӡ��96ぶ�4���~���s����)���1t����Q�t袰�>>��呷�/�/{>�B���s\8��gs؏gR�3m7,�)�F�\��?���i=�5X� �3� ���Ne:
�/�m�Th�4���fN�	����E �/h�nz�{^�7��߿_?�!<����ޥ<j�}����NY�'C��������<Z7��>A��yz+D]����9
������";B�~M�Q>�G-�5��R"��W��7AǦ!����<��}�,��g|��'|�V3���o�i��n_o$~��5��"����ji�ٸI7g���_� W3�`~ۙ��?��B/���Y ��a|�XW�݊T�3��<C@�R�s+mGyD�V+���s��;'#�����{��/����˨F�\RRצv��h�Ǿf�--,�`n�`fR3>�2����A�+47*���՗��Y�L���j�N�,���{A\/������b��}��Z
�&�u�� �ֵ�����1G*)+#���L��X����}<�Urn�͈p�pu,�sy�VXdW�L�p���&�����t/Ĉ<��!�W�41��h�z�tX����	i'i&R��Y����h�>O$n��)ؕ��[3�jg!*��د�/�@�w�G���7�.8���	'U��ї�46��7K~�[��.����ؐeP�f���	����(U׬;����潴����}����4�'<%ic����/R|��K�[�/��2�4�%������t�?�-���֠v��2��ٵ��Ղ�C�yg����Y6l�#خP>��yT���V4�k�y�4g&$5G1��ѷ����d�E��a:� ��?�Xo.�8���9�M�z�D���e��NP�Q���W(�0'>.��į�SJ揮/=91�/tO�E���#GU�J'� zk�A�}�߸|?jz�����z�1GFFf`ż�{��i\��R��Pl:=@D�����k���/�~5u�N����V�T�;���4�=�/?�3>�.Xj4~�ߌ�"�L����	#v�a,zsb}���9���Q�e�JE-���1����u�|_��3�֠����������	�6�$�?I���]��+���|��u{8�����K�T_�(�fM��ҋ2'�d-l*����Χ��WJ���ti���1�<����(jV[G7��m�t����o�(�<��9ڵ�nh�ʏNAn=��ޕA^�Dlu��"�i��F��j�~�3��|ւhKu���(Y	:os�3�5���\؂�$mr~��I��u~N)�ҳ�I=�Z�O�7�R��I)��/���b	�+�M�����xѫ�X�,?����ou���LB��Y ��ݳ<f�8y����L�*�	a�fqY��fh��kUII�'Cǃos���?X��{�"r���\�e��	�sݴ�ŏ[�d2,R<�O�MҒ�������t2F%{'�����Y5Y^\|p��7u�3�鿯rw�� �)�����.�?���,�����DD_�����CR��E��b�w��ق�eZ����Q�Yff&tpxtT�q#�Y�
�M�����s���<�{]�)H�hyK�[=���6�]����y�lyg>��:�|-.<C�%,����t����^��E�I�R���49�,�xd�bO_Bo�e�@Y�@�;J���}^��@�J�i1��^_,F�i���Z�i_c`�Q�`��i�(��參@\k���QZ֩���Li��]�{dx���<ϔ?�%�ޘ�������9�Gd��	b�e�A�s�{���(�NN��{y�(�a~nnGu�g�J�P�����[�)�߆��U����3/MӒ����C�yQ���)0���I�b\˶�*:����KxXB�a%�BJ��NS��V��} �R��j78�(4��`Ek�0���Q��l���{E,�Xv�v�9����[	����u����:~����-�e��V� �5�9G!��:�R�o��l�_OT�:��+����Է?a0�
��b�`���
a�������:�b`Cd�A�L'LQ�E��	9���+Dr��=��[&Vv(i�2�a��rL��6�I�v�}*����V�s���h�S�W��q.�	9
�!�iH�u�wƵ@S6���G"C��#H'�G�U�9\�Z*D�`�:ۯ�z �M��ٝ{�K��RXZ��UzkQt���X�����,�|���K�[��N���cKt���Y��
L��R��A�uO{�k�ʁ����d:O
�9^g��6����0~�}�I��$�����Q��5OvBGQ(I��""'7W�\vF.����xſ��ۡ���&�`��~���~K����?��3�IN^,u�Dz,0��2(�ĩ.if�=��e��F�?.���J:���o��BTkP��}#�lOLa�w�����p�<�	��31''���gW�>��9�4l�6W�PX��_�et�)T]�?.%'P~z�cdd$ݾw��y�s�+��n��6�����Q�9hP3���� �����J��D{ �s�;�A�K���Ax�Ό����{Ή����Z4NCV_귨�%����	���xG[FC�-�����6������"� ��	&�������������U��!��qv~��b�#z�l�����p�n�,;�߹ j40���c�70X}�E��T��vy��+q�t|0��L |�W�/t�� �ݴ�D�20���t��þþ��F������0�#�r��;��F�&��'�����^�]�a��U�H cGb�_�R��]5u��w����#�宓��f�C�|���/��s;�;#���L/?��G������`�/	��8�x�V��%� ���mv~x=�C�$��4bh�b$~�ޜ&Ee��`*���9�B�:�9�^{ˋ��e��V	��&�\(��k�"u'���u~F����꿚/��Ө4w��]�rV����JB��j]F!�����;VW�T݁Հ��!#d���?�����ӢGK�x��l�x�FX�<��i�3�#�yx2pZ�y���P�*p>�w�N5�z>�%CM��GGu���Z���
ݍ}y*��i&*Fw2(�[ֵ95翉{4��\w�w�牊3��z*��ӄ��۔!�$���fuN����ca����lJ����C��+������C�"č*}�Ӏ����������uq��)m�a��/�jg���j]� _����dq;��B�D����J�ˑ�]K�]� ��Bi�D�.�;�����vK��7���>=§��Qc�^�i( 3���5>��1!��m���׏��KU^)B�y�
A�\���.�Q�+���F˳������,Ӏ�`��ո�/_�Q
�J�~�\����Q��]|<`ݯ�a6���3��G��~�$ϔ'_���u	:)�^�Y��x��We<뮾��jE{��>�.���K���5R�Ni�����d/uz�7�=M�'0j6��oE��փ�f�r�؟?K!��`�~�m	OB�N6��/����=���Lu	&�Sz��w	�M�Y+sQ���Q7�b���)��x�$%��<���V\r��po`غ\]���bk�ͱ�Զv6�{�X�ɹF��k��4��t!#�tlw{�enș'/M��JH&@��%o�|�9�1�
�Ha�m򡦦.X�[��8Cgĸ��;�G����4ΘMIB�+��jօ�������te�"�� �ʔj����s e��5C���~�����9h5�x�M�F���>!7T�^��/&�N�e��$�|�q+,��?p8<�__��p�/4Iȁ�82e" �c_����@Y��t@p�$ә2�, ���N�J��YXU�|�4|���B��BÑ�����PV��tr�����,�
�9Q�lY�õ	�6��)���B'f�$�_Pa�4����f��ù�oX�h��[��v��]B�JP� ��"�*CθX}�ꃗ��o��w���٨�^g��B"�6T�;��t>5_���r	 wyΘǿ��%&"0�@�c
k���쫸\~	�<�0���a�'���3����_i�N���o��g�X4(��+�!�YM8���`ζZ?��'YEst���ѕ���9���+�ش��P!���6���EF���H���~M��*�p8tt|��@��^�wh"���tJop�*YN)���4oF��ΰM-���O3�`kF}9B-L:���'BX�5�S2i���}�\L�ŵ���6�2Gկ��}�J��^p�P�A��Q��`�{���*W�v	|��F$v���Ȧ��^���f_��VBk�T-��h�Vq[�0������ ����[z#c@�G�ǽ���d<Vˏ���۷���]G�0�D��*ӎ�/O����:�=sa����%u��(����~:���p�x�
���**�!�
�m��d[��[����'@x�>vW!"���
_�GF;�њ�6��>;w��kw6BP����M^��bXM�p���f��I{8K�KƹW�	9��GvP"`W5��p�p��y�M���+\@=�>a�6����.}�eX���%ӭ���Ac-����/�qo}[�̸�&\zV�Re���f%�k@����^p����E�7��2�M�}�)/B������w��{�>�ӓTh�=�mR��nge&������o������!@��pu'�|�-�w�r"�,6�
���^��{��	{ƨ�/�?[W�*W�*��(�P�:d��?!�� U�p�?��3?*A#$������������5���㓅Z�����]�=l4~�ݔ�/���⮮���ץ��SL��Д����	��<\���%���4Ȩ��`�/v�U��\����~�0���������S���4���W g���eW���G�W���+7ズn.������<�į��-*��rg<_:�:;�L@�����9�`������U:�u�L~�u*N���������x�Q�ή��#^��u}}QΜ�+|��z M�u]w)����9^�� �hɂF
u�G�|||��YlH��P��&֚qßU�UW$���u�=�3�1��h�R����@\{��gʾv��.���D��V���B��W�Q�S]@򟟐�J�G�<��&���6��Fю6 sU� ͣ<�3a�a+ U�E�̴^%%'G��w�h�Y�R�&&&���P� ˂�&���L�uN%�ӳa	��=�=l"^[2�ΣD,ഏ�Kh0��z*.#������DН���8D�Vsue�b���meC<zn��������B }?74�7Л�J}L���1B��H��8tw��o`�V@�����WBэ֛P���v�\�84���#ګ,��*���8R�O�9�{�;P��{��Sl��q���v×�5e#_�(/,"ҭ�fn.��>~� "=�(���X�:5�����4 �)Ӵ�����H��w��nŋ���dʙ��}�E��Jko��Zr	��$ ��Bm�����e��NC.���v��I���ț������W2|��n�,��������%�UPm�< ��K���r�j���[�Yʏ ] �vwיv��,���I���I�i�O�|�j<��^1�Ku�A��.s7�̌�q��$&nT��8R��b9 �	�:;%�vQ��i�o�T#�9
Z!Ǵ�ܲ>��%έ�o<;�����f�8iy�W���ᖂ���T�T�f��+Q�U*�����t�:@�#���W!�Ζ���X;��-����:��hHd���k�3��S��N�ﴂ��*�ȿl
�Z�r�G;����q3��������������o��v>Eu�x7ǚe��}m)��E3�9Ң��ͯ�Q������ps��?6�>PfVJ�������X3nO*а�r�CM�5�zB$,tsk&��'��8����G8���*uh�_ٺ�&����}�6m|�Y߃*tQ�{�Nrv�"�3�!%#���)�I����6�.�,Q�&^�-������̙��Xe���lk��==k	))#����K���m�SD�q���՞omgg�k�No�:�@�˂%e}��->|	��i_Ӎ�С��6��H��о�|$�8M\MA[����x��G��@��E}T�-�Nq �w�3F���<K������)1^��A5='~dA���2o��&��ع$is��<|F$911a��k�B��c�T����!�JHDD��0����d�z�/>��%���$F�k؀�� �+?x�m��ۂ�x}��{�tW���j�C�Ru��/��?�!������x�B@� �����mZF��j�&���S5j�X"����Hڻ�^6Ϻ�������$g����at�i��}�UTF�(� �@��`��]�q;U����B��{�����i����ǖ���{�Q_̣x�߬��>e�*'���΁�ׯ�?���fK�ק�
���GE[f����$������J@'#t��OKLhDj�Ԙ��XxS�ax'R����Bw ��w5hF��=&��ݬ !	��5er�	�H���>�H�2��\�\��	,Oη�9ǁ�+��~�8�DT�T����]N��p�+d-z���P��)�;�GNNN>�4�];�c7��O�������6B�B�|���Ϝ?�bl��L���g֏��R���^9M��Q��I�uKV�o�+	�2����u�����E�U�udј\yg=�Z�k�l���pS����[�l��,��i���_�������Ϙ	Q��
�����<��|�4�S�׏.q/.-��a�I��5�R^�09�	

rX����mf��=����-6.~��:[�GM��n�.dV:���談6^(_�A�7w؛��7��%��V~�P�э|��a\2��M�M�v-�WՖS;{�GM�-	U��0�Ǐ�S��n޼	��kr��>���ܕ�o�����|��nC����q^-�x��?�F B�-��ݰ�.�,dH�+J!-#C�r0鵞o�)R.ho��1��(Ǚ�D��	q���s7/�=X�pf���Y�CE��g_�n������j"w	f�-��|r���,�}wL��O�6.Tn"�|�J��ի��_��Lk/
nŽ�����ucœ���xz� ��tu ��|{5��],���[�SL�Q�,��R��*�z�m���w�E����m
9������O�H@5���� ��&
�K��eX9_� �-
$t�I����]Y��5�MP�
�E=��{�n�8��Y�C�^���ww�e4��bz�'��%�+�`ħv<)���eW����=�g��ym�>)��$����faa�{����Z{���p����.���/vTX�* �m�����ָ�\�M��>'�eJz::y��@�Px���/.��$�>���t1%��k�9X�J�H�Z?�+��^9�{� Z.F�J1^юS�V�������?br��3���b����ZՇX]�GF�BG�᫈Ɗ�e�v=����9S^U��G	�D����1������f$.�L�G��,]LO__n�]&����\,\p0[KYc�����;�k�a�U��egg2[)����w4BK[Z��x�:�\�ة�_9�V&�Wz�� �?e#�ۼ�W�}���dffV�Y�A���1�$�eg ����s������;䷉�)�2>�O������L	)�We��ލ_�~o}z9K*5�2����>%f{���Û�C��C�:�89t�99i�x�j|Β+��
 &��^��s|T�7�sX��ܷtt�䫕,W�,����) l�t�X&S��:f�������>����{3v�5�:* �l; �y�) S�����$ԃ���2�����u����T�j\Y�r>�n8���N`��Gj�K��v����~#?~|R˿u⬣ma�p���8��!�4F' �n��}�T�1.�L+��o�aWLED����Ǯځ�		I�zh������+b��{/b'ȚڟK+�:\�Pܐ߃�B�c\��K�Q0�~�(��a�5f[�IG��2"��knm4�l�K�5&�b_kO���j�ʁGӊzj\@\b�������8B-�����~0����sg�pZ��_߰���IM�
�m��v���"\d��!��2�*Bv����lb'��4���0�[�z�/m���]�q��|S ����MB<�m���+<�w�������ٶ�`��n u��l��ӿ ��!7��q#`�ç-��w��;�g�G'��B�V>ՠ
ɯ]����rB�33�Q�!�]��7���-�{{	).�^ϙ��{�o�q <� �İiC��|��<h�~q��)��]��lx�?���Y��2sD��A�e�Zy4Q��@D�R:���d�z-r��|��̎ҟ:U�(�}��<�>vs3M�p�#/��sKˎ]=�b�2�a�����V������gcu��zU�fvĝ�!��� ��k��Ŝ	���_2�X��[oF�4��e���W�{�5��ƨ�?2���7��dY��K�\�U�?	��WW+�=ob�4�M�� ���N�i�e�g�#��z�U�D�%�2dXO��l4�pl7qSP��j����֭�o�p�R���zR6f_l �ӫ����� ���pO��]�T��8��#�"��j�q�'G�f��+8�u�ʘ�ړF��0aaaK^�J�d��TSid�p���޾���SzZ�M�$�j8����Hz�b�+Ā�x����k�����hxbb��.j5��Ғ�SU�UĿ��`X5��oߤjL �U�}����N�$d��u�aMfM;ꂫ���"��T�w\Q@zG�J/�C��"������^B���C@D�I	�tBB����~�%?�}w�9���}�s��H�UKo&�e�Ϟl�}���l& $T����e�TY��������9�Qd�̯�GTp����(C�\:���Qz�q��\�cy���ّ;����ؼ�����%��	:,|��'��CoK�)��pD�j|�#J���jq�:���[gQ�_\RRQ\www�&����2~E��^]`��!i�����2Gޓ�f���$�g啕�_�̅�ea�����a���_ �XI��]�u.�^V��[�o�QÄn"�I�}��N�1�� 7�Ã��l����nTʲ1�%�j���Y$0z��_#\�cC#��H���eM(M�0����zJX5�w��s�'L��ҏ����4�D0���p�Q��@l'	H���R�ԢJ��o��q�0*+ݒ2�!i�$ͼ���t���/D �Rew�.�+�>(�����'��t?;���\�����E��z��bf�߹�08j3v����� �CxWb\gIH%�{y��N�XD�o_�~�<}�9�{������kc�9p ��N�$�J�sC �4;;`��,��q&{����z�<]䔑����;�����t�E�Y���P�SE��ڽ�ܞƋ���,��O��ݝj%�j��:C 5��p���7�VҠ�L�a�&&S����j�T'n͜{�\�����hZHXg~f��hg{{�����I�f۠^��h�-��`I�LC�s�� n-d߄��T���]pdI�|\��N�&/`���_~<���~o[��ۊ
>|�sV�E�w�τ�uL�?}M�Do��:���D�9�������ꇠ���I�����|
�K`2{��N!�@����;�T:��..�����Md��y"�G>跷�2�ʋ�+볲��%j����c(�1W9���>���������p�����vN��Q�h�����67���0���Oa|#Y߆XܥV�3�4wE?��;�QMoo��^G�pIn�_�*X��;T� ��A7����
� �C��"���3g/.�d�Ũ�� �87��ep�b�&���r�^����/kNtWF������rkRcufZ��c}���[�+�g;⅄�r �Vxs�Hw��P�\7q�o#�jܳ3�V4�F��6sA)��bêvA�*�b#�&V�����e�D�4�"}Sά�_4:F۴s�j�d[ĝ/������>4My}wf���9��4��Ѩ�����c߾D}����xM����Pa��-at@�gyJ�\8G߂��1�o:�v������u��|��/Guս�S�$�aĒ���b��B�ޞ�~�p��p�J���;]]]�׽K�|fq�~�b�Ĭ�D�N=y�~R@��{
�H)%%��� �wG ky�HɌ�õg+9�"?߮�ʂ�˘:DY��#�a*O�Id|v�Ī�q>r�U^�Y}zNEU� /O��<Z����k��p�L*_܇�![�����i�I 	�a�gΎ��4�0 A֛�Q�WI�-qƾ�&��w!�8����5~D�4�*[�NS�)r����z�Ɗm��g�aLӑ4\��;���N+s�� f&&'������G�^jz�.+����mY.dGgu���!��Ë��o@�r���Yn�^�}��_�v��U��$K:C<��nZ7�ҴP�g����\�Ipț����-$h������� ZS�W��oit6�9��4���;X�N��ϷsrR�R�])���\M��a,��c�eQ��9pt��p�k&%w��yڽ��謫���ۜ	5eX�߄cll�r���AqBJ� ԥ$��*D#��?�u	@�(c�I�J��e�����S��q�5�{B	-EA���'��G�l�O�=mH��U��G�K>���a��@`u~�n����\-�k{�o[�4;��fu=?k����l'|7T���Π�����Tϟ�f7���2n��˵0kkP�'��2���&�`��uP|�Sv�a�`��]�3u,�ք�@��\�� ��2t�w-l�lncn���d��4?p�Ls�C��s�!YK�ok�WC~���Csq���g������`f�郌4ws��EX'»L��ߒV�n�C�)XE(�)����e��nU<����n���ɯ�$�-���UiUQ&h@�o<�B�eEmzU��JRB���`	7�N�_;Xa��8˲�#�1X�]��LP��z�/���e�r�I:��Xݗ�qPe(+y5j��-q��]���Ď�Y�d�G���
��56M��}�g�pU��B1t��&M���O��t��e��/0X��\�:�!�"&,-(�8g�j�V '?�u;�����+�1�݁������i(��w��V���u�G�,�+�#������Α��ϑtk���j�)))��46F�cu�ɇ^��݅��1_=�������5_)��p�]���7`���V.���dv�޷�P�(]�}J���IIZ����i6a��. �����*�������a �����������%��ס|,��ϖ�ĄI��������e�>��	�i����ЪR���4|�h��
�ņ�}/�z��@�P���4����!�Xd1`Кyʩ���pY,!h$�����A�w��Vby'�U����g�{L.y�����H"4�%�����ydVV�����-�<��:C(bG,�ߣt��4$R�jj��C�(��Ih*�Χ�����\��bKb;��B\o����q����8�$�p�Mi�Aԋ�Bac=Ϋ9}6�m�7���["��2c�.\\\#�pC"E�6�=)���~����+p��kY�����<��@V���["�uj���R�V̉�x���+.4�vd�-���5��L=n^"B����GFB�� ڌ��54�T����<"�`����⧅z����?��W�SN�<i����Q�xr�D���>E�Gj:��Q��l��ɭ~-�rhI��L����N;�A�ѳ��8}������h�{u�gaN���A`ͳ�J��ޗ�TƵh��i��X�(�#�s�E�-CwP_u\�1�YTz�Mq<����/��n���>A��p̈́�;�++g;�(w��Gி��ϧ}����Bj�Wb�3w�}Ԡ�Y6!����mK��
���1�(:�3��J�b���t��b���3��XIUG�������~lnV���`�wQ�B�if]�h�~/���D�i̴��f��>�Ӌ�`˄
�|Sw2V�����x�Ӗ�F	]}iV�ۿ�X]xS�g/�<˚��nM�
3Bl�`�w	����
5Y}�h�sX��8@��P=��׍�v@ެ	�8,i߾�H�=^s;%����k
�}�Tu!\jw��%���0��u�]g�d���	`9W�w5�NzgQE���Ź�$C���N7��rz�BmH��q'zdS[��i�
����q''i�G9�����<��ı�\.eN�r��X�W�V�.i|Em�#���c�ӵ9��^��)�)��[��V�� �rP*�Ø� _����"��^���lo8(���K�����6�f������/�2|���D~��>�Xw�/�8üߟe�p���=�*�%(-�����궐 �V�,��bF��`�GDK�ߧ�jN�����>��l���åB���1�u���6�6!/ �_�gB	�\�3����źBbbP.?`ٌ Tmh�d�"z�F�3����ln�i����o2��'l����߯=&�ӧ������2(��.
}%L�<��u�a7�n���y��ꆧ$b#X�
�ߚ����<���([�<�+�s�������s��_�h�Tt�D�K����*���*���@�	�6���R���k��O�D����C���J��l��:<\�\e3ۑe�AX��Zf
��93sss�q0N����"�	Y�U����7��i�W)�������0Tj�D  py~�#����G<�ħ��e7�m��{k-�|2l�,�`�Y۴�zTqLk�p�G(�$���4n��3(w�E�5�}��ٚ���q	����MC�0F��Z�ow��A�۴@3��QZ��	d�=�FE]z���v�=w�� �رmB�Y9y���P=_&�j�P�������*s��W%S��R���uwG[�}5J���� �ѣ4� ��v8��� ɺ����\d����Uw����GeJ� �(h����TNS��R��%��Z����A14<�J�ރ�K�>��vZ7�S�}im�g���o�ӣoxE�z(/Dz��#���ɸ�������Z�J���?v"j��(��,�*�<�τ�R�7I�v�1�>:BͩJy�m�.�vԿp��[%���AC�Ž�4=@��_w���X��W�$��ckҀg��c����ts�?�RT�q�lT~?��p*=���w	�x��R�s������e�U'�@�]ϴ��$�"��[#���w^��<�ӀQ*��bXz}��ߍR�⢢��W�N�Q+�b���q`8�}�p.����[" �(��f4L}��\�]��U���M"8 �w��m�֥�:^��k�F7�)�+m�ėo���Ti7K�*2A������~�#9996$�ٿ~��'�P[�s+��;1OS��ۃ[S���f�R���(�����| a���]p0��^�Sк��!���4�cM�Z��Kn����F�x�+�a_��IM������\�?#c��#++�_f�vE�����:���x��ZE��.��J�b��DSW	@영��w�Y�S�u��Dg��r2m��au��������Ss�l����͜��,�М|?��QSV��	G�e��[.��J�+ԓ����A��}1�Y25\�+VxS�07���a)\d\���Y"��.g,T�ݔ ͍�YY\D֙���ct����v��^��x
�,�#���xϱs�OO@����ۖ[��{�5�-;G�����E�i��G�#[�  ���y+�Ń[h ����6glE����z,��N�_%��������퇁>u���-z/3��sgEչ-FC|�eУ�U�顱��@KA��g{ٹHs�t���Q8��61t�6ko$�rZ�3� j\�g�V�Xa�$��@����w��t�w�UǊ�����Tˍ*� D ��}s�]w��r�G�F��Y$�*����0#w4XL���D��.�X_��3�j.��d�lE�{����f�O��hll����-pf�:��H.�fl5��8U�����,sG?N۠fɃ
�(�����ClGױ$�^x���؏-���;���f?��g-�OKJ�r���nm��H���i�[ڜ�vV��ꜱ�2B��F}0޾)����ǁ>I����|��r��ˋ��%N�ܥ��|����VP��1Jl���V2�-� #޵,M��օsk��$��1�)��r*],!������	ɳ��Ϝ9s�2hVF�D�ߑ~Pp��Xe�i��]�ez� ͓�^���xs���� ���pW󕖖�D�KNA�;������g¶���%^�&�?��M������w7E���\��  +ц>*b,"�#��\��Ãj�3�Y��c[.�b�b��?��������v�wĪJ�&K�j��F�'�$��TJf�6���c=��&�kO�.������#�<�Ӛ��������+��n�����.'��O\�������muDĈ���!�5�R q�D"�
}�[�`�~F:Hm��Q��T󶠧�Q�,����WF��c*J\�ۈRk�b��z� #�5��YjM�̃�ڞ������4����I�X7ť�$[l[qҞ����cb�*V��\UĔ/��u���RQ�'�eE�}�����˥�q�Ôp�l���&��G�V�ǲ�v��_|�˭��>5����ig�i��r���@A��6��	*N�k�+O��t��%5k�Pv:���"17..�m��H>��-,���M������9�?��/�병:���e�,�Q	]�I��k'*�,������"�1��/K��	+xLɄ�� �7����m�W��8���^�mm|���������x��P��q��� ]��|iU.���?3����=QNb��&U��H���6�J�Ӂ�3F���xxx;E&��bw�:o�#I��'�o/|�0}�/����NC`��nٛ�D����\�LǸ����'
�1[obTbq�;�{[���΍b����x!\ _�hl�tE�h��:��ٌ�<��P����7�gM�@�2�S�p�Umŉ�]$"�^��ޜ�����l@&+**�	vn�����饥�h6s��~}���?z"�b�4��2{12�7/�|������E�3�=ҳ���B��a�i���w,�(-��7�/����L�`�kz�{x��##KvZ���da鋬<<t�>���ަן��h�.-@�:�~*�ʺ�o}�D����*�rz�k�}{�y��S�*b�"��HU��I��W���I�*��K�p�ƀ	���n���_hg J�仨I�}*�#�����4ռض�m���⼴����
��ws�r��5��d2�� �۬�?�c�ҕ.��L�X�)I��&�:>^��&��}+j�vd�L����Alŭܖc=NWFO�#;��	 r�q+k�0�^E���2��G��񟐜�����X���l�;��κ�4������W�|��'����lB�#���.��1-wH�Mէo�˄<Ѐ�N��!`�W��NU�m���%�F/[&�BA���m��Qk Y�>�彄���HV���k��(+`��-��3"�������`K]P$��Ь����D�ؑ��10���iZ��j�">@L�&�J.�����C#��{����;��ڼ|�yP*���{����"�	��%�Xׇ�!�e��)���k����*���أm�~��������V��D��Ϭ�N5C��wv��3L1K�_��x�{UW��S�ȸg ������5�?��ɘ����#��\�z��-�I����=�@jA�����É%;L�������)UI1|K�����}�9C`�~&%(�0�.�
�ٚd�ܚ�)Y
T��~��0�"^a�>�XŜ��@�%�>Q"�J�B��DL��ԙF����|$���P�Z@���76������)��N��&��	n�Q~*��￙�j�����|�)�Չ^i����:3YenJ��twFv��8C������r�`���`#A�u��#��/��J6��A==!A�l�Cx-���\�i�[0� ֥�hv�j�'��x��ㅟj�>�9�rb#�&'���Kd���K�=��O%[�A�Е6�5V�͡&��Z4$�i�ո�l�ގ�+W��-\sDq�}�u�p�0��V	�co�Yvs��m��5�%ٸ���I��0r�D�?�����b�9���Y�� ��bccC�u�w�˷�������TF2��1m����B����ݐ��{4�ׅ��">�H��p��N{{{붡ܯa"�L%⬼��k�J,����~�1$����^Q���WӏQ?Oq��n1��'IڷI��o��v{ۧ>�h����鵒ޠ'��E+A�#}$���o�����߈����:}pC�}ˉKVە��9-�裴9�'}�1	>?l��V��H�YHٰ��1�S@`fo�}�pQ\|<�䀔�hl�TxE��;}x(;�B�O$��L�%�?6�P__Lʓvbz~���H��	��0�%�j�.���`��7��G���1�|�����"��$���)����1�b��������9�s	�o
�
��k��?�Eyy�!��J�|���ٟEl�r^����x�sd,�n�(ieeu��;s��yI�T�⦪��>�۾5q����j�$����_)�R��bMդ�>�\��;��9^N�Dz�2;�[�:~:��}�����&  ��|6j��{�5|��>�dlYq�4���_%�Oݕ�Bg�o��́�S`�<K�D�m̻O}����jxX_�36�.��o��q>1)�=yO�S{��4��I��SZ�*��)@)wJ�rfOn]�;�g������)ԁ�q<���@K�$~�O���?M���|D�0R>�!?5	��Q�%j����Zg��{��<�\�[P#jq�-amN���U���56�?%F5/}�( l�я=����D��	���`o{n_��0J�s�|熹�IZZZ��,J1'3�b"�������� Q��r��g�K�Q�~�RLO�TW��)K�z��&\��@o\����U9�|6�+�V����ݲ��d` ̊�(< w�D�W��t�G��]Z#
#���ЃT�w��_i����Q��Lz~<���J�=ҵP��'�����/_H� �]�7Tj���2V�S��L���s��a|Y�ֳ���VhL�uZ�B}���s����&{�#�^��D��`�5E��\����Tsyx�M�.I�|1�s��G�*R�ȸ�bWlm��������&�j�z���44\ש
�q���,@����ј���VsW3��V�ޭ&W/�X?5��0���,%&��(���w�h���)�M}S��|���;0�C룚��p���ٰ�����{����K�+�z6.g_	�HJ�N��)sL�0��~�8������=�O��i�,�?���988趷n���AxD���|����j�������ǎsչ�|�)$��B}{Y�dK����6'|�a��(��b���	j'�a�;U���ջL'z��M�yRP�+�l��Q���$�S��lu�vP��r?�G��#v(�},ܡ5�9��O�U��MA�
#Jg�b7��Q~I�`���IHe�TS^>�Į.����ܽ�c8����nc�@<��L��ڇ])�Yx֟ߴ��V�W�\s�+J�:b��vq`�d-���
�_{��rt,pK��jqq147Rq3k�ZS��$cAN|#���~�|C���#f��n��/����SE������VHI����/�2X�菝%{t�Z��L�1c���4�_��vF��i\�s�����E��Y�͐����
���\xډh/�$K�U���iERu���S�9�o�J����vNjy}Е���\��ܐ�"h��$�yuQ&����6�1w�j|���>�i���2L��7t����^2��5X��i�k���<]��E<��$^�,���Dj��o�d��?�Xt�����%������[�$�t�X^^�]�����:�{P���(�N��>��#j#��I����V��G�½��e�Bd3 N�=΋8�p�j��z��Q��iaa�;�ș�L��}?���4��T֯s��t'�A.�k��������҇��p�=D&'2�����Ya(��S��b=������F�7���o�KF�M {{^�	��)����y�t��g���{Wk�>.��@,<�l��Z �4��f�*X�&�P�9������4�C��z��\}�wNT�S��<L9N���
����ӡ�I��y�Ax��újb���.�E��J�}q��e3fek<+�{-#:��H{yq@����Vyћ���KK�A���`�6��',��� o��G�KXGlw\Y��4�7���yw����% ̎ﰀ���|MJ�}����\�H�؟Y����l���I��a�栺c��J¯^��g�|���h���L��p,�S�v{���q�ē7hA��
<lm�R�H��wa}�c�l�b��VAn^��+�}��Տ�qk�;��V��X�
`D����:���������BrVS#��;B�L�i�  �9(�:��Gl1����T������;(h�f�����	I
�u�����}�m�~~=؃t�:O��i��&��&�bkq�D����hԪ�˟�.�%�����8֪W�s��A��+T�K᥅�[���FY ��w�F�k቎C�o�IL��U ~"��S�D��wu����T�ء�^��1W@��#3�]$9�T��s�1F䇸���m���.��F���.\w��P�������1`�L��t��'��"k*m���pY�ć8�����U��0��6��=�;�]]]���$3��i)�����y�8��=vdh�q	��xI�cG�&/E�E@^������t���0;�r_1Ҧ�	�Q���ϟ/ǲ�&IL��oM�{
��L��u�7���:�+�[(���ZE��DE�W4�(��'�5�{w��}����`���:�A�`M�΢��>@U�W�G7��"�3�0|\�e	Px���gk6��5���`I+�2�~Ocg�M1+����EW���E �����ee��4���,�c�AAA��j�ƈ{��i�$O����|(�y�n�bbZz��B��Yk���{�e�w�������<ǓJK^�VK&�`�1�S�|{�Y2�Y�(�c��mV��4@p<?�֖�B�F%����cv_�!�iLP����W���$ɂ-|gML���J8T/N],�M�d7�975t��|W�<AqP�d�����,f{�n�Ch�=�W�_	�[#�^�����x��ڀ�;K&�І��胣mj�!qw����'~�dwc�7z�A��ބ��t?��	�M����@��T���y�M�����FZ����i,�����(�p �����
�`�C��'�_|(X-���uh,��Z'�?�ځ�L~t�W��o����P���)�qO��I+�(�ơ���֥�ܒ���~�����lУ�����V��+�ż�8����	2q�)�Ѣt.eQ��#gqq�y��Kz�Y�= �P�6�-��5�x��OPk�����R�>�?�X �ޚ3����*�I��h\ N��Y�������ej,UY��Ej̆�aް�?tZn��k�^����{~�Z�$�P	�'���}�f15`�j�ܯ6�!wI�,L����&ͭE@H��=B�g��3�w���[�ߏ\���I��M6
����{�H�}ë,��r
	�:�m����% �Vi�\��1m� 饤���"��1�r ��y��Y��QFzlll�VD1M��\?zT�K�������H���)���iʈ�(;h `�Pҋ���
ƹywd$Q����mO̗N�z�y�u��2�V�x��?�\��m�����װ�s��Idq��;�X�֩8+>0�u��uը��Y1����p�U���-��
�C�8��j*�j�<#��V.���_���A��i����p��~��LC��6 0O}Y��z�}*/	s�4���;�q��I�wj,�4�g7��#I[��~�4�p�c2U�������g:7hH���c��<��׭5J�:��܎�}�}k�B4�Z��N��CXX�=�8�0w=1��P:MP���Ly$Ǖ�_H�v�at��g3�|3B3}� 3nu�v����ş�n���c�����z�e�6|�E���:��q�i�������I�=�ܳ�M�?L�ݥ�4�nB����������ا�O�_4�M#כ_?���tni�I����LȄ^Y�����3s�	$�;�����̮���m9c�^}�+�����!��̏%!�`����c�@��iٷD_�k^c&l�������P�i����*`2{���!%Em���Ƿ�K��S��UO�?��^�";�����H��AB�ev� "Cw:���\���q��<�_hq���C<9o�oU�0�W/Mq���>�HϏ����B�8Xǲ๗���cθ��2���߷�Ӑ�8 ����;�.\�RVQ(r��y��-HpW#U=8�N��a�W͛�Rw,�_��NM��`��@.�����<�SK����7a���BW�l3bM]P� ��ʇ����H*�9:+��j�nma�������ќ#9�a#e���V!�HVh ��l�)��I�u�<3�h�欞��Z"�rGxz���zM��}��e�w��Ɏj��qq[����D�C�2�� CuO�Yw��=�;}�T�R��fT'M�7r0�ڍ"p��^+�O����܊�� ��ݐ1>�z=R �?�K�����(9��������~�=�� ���Z��Z58|)1ދ=�:֝�N3�y��D9B�h���K�6t��ebT�?Mw,�l��JH?ށJV�q�^g_¾
_�QW%ïW9A_�=��9���Gr��⏜ZB�q���9�)�t�q�F���:�z��]d�� _f<���xd�L���>9��a�Dg�u����9��CVV���
v���i��X���SfC��U��a�q��Q��vp'q{�\�%����`�Զkm�`�����V������,bGY+?�-Z)3�3�^�(�
To}�W���No�x-=�x! ����|P̓ӄ�H̍n����;�`����:R��9��=e՗�o��q2�܅��𧱛e�	:J{���+�Q�z�i�)G���!���Tx���v8h$;����_�ulz#m���`|v�M�B�v�d�_��w��f3�P>ii[�1�M��'���.<R,�����;8���H%�v��<���Je&��1;��Q0r@��eH��T�sZ�-0��s
��v�r�fOʾ'��C#�ʭ�Gj�$�(s@u�~KZi.��e܅�^!�f�,�W)fV�c�V���:\�a�	A�+j��G}/0��m���x���u�,���`��J�4����c�������=m���
سV�S����=�\N(M~Rom�4Ec{h �`��x��"�6�Ǥ��	v����z0O�Ȇ>xꑦ`�
wb����]�A�w"�}q���[����f:�O�o/��3>�;'G�<�ä��z�T��5��h��L���I���e�e��>�����}�����di����2�w~��/ѰA6��~�����]�!S� �������&�q��ٓ��	B5�_[[�c��N�DPa�)Mǳ�v�Q&���D�_Fp��i��$SRR)��b�yz4�J��J�(��@�f�*C���D��6w�;\{{�Q�zV���(pG!x�d��E��o�4m����>�}B�1�=<16�.�Df���#&���vRVd��h?��b{��Q*��n����C����¡��������[��N˝a�h�T6��/"5���5
�geE
������ж���~~���&*J��~W+�Ϳ��$��KѰJ�l�����9��$��ZwBr��<�����HZ�s0�G$ �p9��#"�?��� ���&+��Hl�c��G��b
±��b��Ɛ������� k�4t�����Sw�i|G�um�W-15�S��G��Bܜ
Ǵ���	�j�X���,�r��j���� �*�@���jCi���n@uo�v��"���~\	�ng߶���B�ڈs-`U��oa�18?9�܏9�W���̱�;� o����[���n�B�nV]MM����^��l�����klJ��i���3�h7��n��3��Ʒ"#��r�2еUw���z��Sl���}�'�(�<�d�j��3�{NV�p�hhdȳx=���>��zr�R������VHM&`ݣ�N�Ed�?� ��&ѥf��2,7���]U������b��	���T�%�]̷_ɕ�;�?-C6�f����u��WV�9���؜�1�{7Xk�*>,�~Q���$aq�j�\�Z���:��s��)�����X~ԯD)�k�	�-V �r�T{�4t��C��%H@X8�M������"~Qz�'C�����S�I��e��|�=�_��޶NCy�FA�b�r˗>O�e��,z�D?Eף��'L�6��C����ق��$OҐ�!V���m.��@w�G�~���B�C\��C�#,�@�LPZ����0�v�T���R�P�PճR숵�raf���{�5�e�m�u���,��`x�]�P�A�i��E5��4,ߟ	(Wq�J/=��~4m]�U.J�1�+���g.�.���**M0Z�u>�s�$՜{���v��Q|�S#��پ$L�V��"��*�q��4�c^(��~' �N��#��8�*`
���<6�|���p��n�+��7`v�>4���0����Ό��d2��lÜ1�y3{��Wc ���O����JG7��/���ן֝�BbG��a-/ŝ>��gl8��'u�N	4����~��YGYA���WQ	���H�����'��?�C�9���M�ָ+����r�,Y�n��'s�,c���;���Ii����P�R��������$/��N�>��Þ��h��b�\Jܸ>�l�?S���(hl{U�qR:$���ׄ�����/ߟ��]~.�o�u�Y��"�#m4��ۿ�JJ[�nG�;���^�HC��u��~E���?�?2��,G�$i��bnͳ²31���s1]��<��hV'Ʃٴ�1�l͙bH�;j��t���B�m�_���Z�q�O��1�����;׌9!I���Z�"%4��M�Q���m.K��>?UvJkm����9�#v�agc��[�IWCC�k[�޳z���[>���1#��xƥ�Z�2w��J�kb�Vv;����.��rxD�l��`��ዚ1�\�3OA�ZZZ���<�I�=�Ex6;%� ��娞�h�8[��+��%�
�����;s;��|n>Y�� *�VMu֚��p��8ދ_�I�7�!{ qw0���SڥN_s�I��;�����阎��w��i��g.*"ۮ����]ŏ��Ȭ,Y˺�]rv�AlU��������w	�o�d��׉*:��bM��ݡ��k<�A��U���e�j,�z�t�3M&�����Z���ߋT�N�ɲ�b��W$�RW�%?��ԼH@���|�A�Gh���py���������D
��]"˫�ulZr+���H�s�T��1�ϥ8OrM�7��%�'�5:���^�R�!�@�����{f��2�����£b��Q�2�ؙ$ҽx���g��)^�ڷ�oy-���+����Í��}�ظ��2����$9yx�cBk�p<=����m2�zp��Q4�
��}�ݲ}�Mv��o��$��;H�޺����i�W��S�����T��_���ꣁĝ���`yi�f��cONs�����Q��snL/����ͫǟ<�Os� r i���훂�������4j�e;�U���tл���ɋ�#h.�Nc���:��"�axdda]��:���n���4�uZ�V��8�"o���$4�䓡���r��KI�x��_|�{��8�aw͔S�%u����S@��@yh��a�}�?��܆�z�F������;g�8�;�b�5�� ��psn<���Yr4;�U
ܑ���g{��Wq�֨�����)_|Gl9j�FǷ�K�+�]~�|[�L��p�ߴ��ڲ(�������}��.���ut؟z�!�I��-A�	�9ո\�碣]���Y[snyYJ�<����W�a;�*��\�@/��Ų$����yO��@�O��hh��Ԍ.�<x�=���@����I�Ʌ�P��4�i����/�?�; �of/�~����³���xGkg<<#b���caa![�bE�˫�vw�hM�Լ�s���ҡ����-���R�q�C��1�3k2��@,��� ڪ�2s�=L�5�\������s��(�D�	��n��W��]��n�r#E�M}���7��ݢgԌ��:��
E)�����ɦ@���j�������Uꂀ�*,q����2S|�>y1,��Z��S�F�S"�c�4?t�\(����s�%|�S���o��e�9{Ѽ� �^�y���˧��n$(/m.�As�S}Hb~�}iq�,u��������V6Z��ܳ�k�xf�mK��aWeh�����wu�wR�If��P�Y�Y����0h\����Qw�$*���)ҰA�]c�0��%��"#��F�k�8?8%�����3�����d=����j$ԔʥRO_?A\Bb`` �Er������f&_)�L!�=��hydYHn���~�M����L�ؠ,�H%����t`�?Xb�Uu��� �ao���*��;`K�!҅�g�2��'s�sVK�r�dC[�!���V� ں�V�Z�K�H]VV����2n�K�ݵi�H|G���4[�ᶻ���oc#���>52�51GOE�kfh���2G����޿�l^u�6�ר�����I���Z��ighJ輻�5�M�;���:�Ö�g�C�vt���GJ�l�� NN�(�<��+Iv;[oΏT`������ʢ�Q5����؞d�[-9.6�\�Q���Zφ�<��������}A�����=�B?R
V]��5 � � ._U��fݧ?v�)�뀫�bԝ�216�y��A�5��ţU*$n�gn�`�����իW��� �L�R]s������4��S������^�e�z��PC���?��x��Ĭ�W�����@֧t��d��������!]	7ln�`>{vhE&r����\�c��'��8�"���xp����&$FF���K��=Е���lii�T�*��H1z��D"ָ��F�:�QW����iȹ��GETz$�X.t�l�Տ�;>�g��+��{[�m��2��A�ZZ1}G@�e���YL�p\�* �H����׿U�1��\�^���*��׏*ZV+k��/^�---}�"`���kL�4[:M��QƝ7}�����َx5����<'R���r$'���Gs����L���Օ���L�S�!S���v�_�C����ٽ���k��me����6NN�GGGׯ����y{{;���;���$��±�[�� ��a#���J��o�Xo@��Wz��**7�o��~*(,tݏL阅���>5�,f��#!���߱(��\6�"��J�3נ֦�;�X���Q.������hGG'''�S|�#"�/��P�-��h����j�c�S#��6'I��"���Յ��KE�Y��E�#]���3ϻ\u蛡� ��F���G�����������9����@��N{�Lm#���5O�_M���ڊ���o�z+��y|�<e���G,,����n\��zf������T{�6��� �o�����j��*oP�f��N�3��LÚlG'p=11���1�=��W�͙�4�a��Q.���_����P0z�{O�'f\_����
��:���\aG��K�+V6�8/�����;/}��S��N�ٙ��?X{�e���,t�g�{��"�M3 +�TT3w�S�B��-K4�@��Tn���o.�Z��	 Y]��,�I�טE\�������w�xoWd�5���s���㯞�����7Z��"�>��jGˠ~�u0Ah�k�<|�^.T}&�99O���틞���bb+c����G7�O�%^I������@A?
�/����L���7�$Q�GhM�Bگ9F�]��PhVͻ}��i
���m���1;~�������6�c����:N�=�Ј��� *
J�����}o�EU���JǉTp&��ǘ�0X#<)�}�d D:�x~��u��	 ������T[ϼ������6�BXR�;N�${�ul5�2����<���Y5Z�����Lb߉%�9ɩ�I�n7k�j����sI�+����'}�BDi�q����� �z���aRBZJD�D@Z��F)�Mw���l����DE@$6!nR�- �����|��k�sTp3�ֽ�{�̚ƽΩ6���
Q���v������Y`4������`�}h8�vw˵���y�b�����!�A��d�d�IQΝ�w�W��<�QG�rEp-ź�eIA�w�����Q���%��-����E��v2��;)��@h����/��%jY6Z�X�SW����Z��#GI���	��k��Q�v�9j��z���w�T?�W���qE٧�W�VW�n�@�F��<�)�(EI.b�S��f�A���k%[�"T����u��	������C�\�5�P��,!
�$����ö�|&���R�>��m�E�+�&S�ʕ��ҷۘ�	�2�<�dx��gp�R��oVW_�a(�a�䗾>6^��y��D!|�!�]��iC�'��f�5U
�6X��좏����Rj�q3s�����;Wάx�%Oj�2x�S�M6��������K1ҟ�73�j� �[�'�����tM�"*TZv�K� �m 8���\R����5j�(r���A.��MjР�eM_w�v�*y�p�\��"c���M�5�����g��+,++S�=�O�S�1��T��d��]Ac9Ӏ)d99�_>݋ �d��$�0GX|J�%��f�kuI�R���s��op�ۼ�6�֝�1��Kb��갦553����˪�U+���ګ];��hZA�����^(K ��r���E���2����X�^k�}��WcQ;�)w=�P�:��J�!�u�3�fNR��.�vnߍ��}Ĩ��#^��=����Էc.�!��X���)�و�n����u��+vŬ�hڝ�R3$��G��Yӥ��6�����Ư�����g��v��8͊��Zo?�a��*D
�B�+�*T�z�EĲc;�R^n?U�`͔�h��@�kG�$q�ɓ��N ��K�@��Y��<��@��ڐ��-�I�a�r����s�s"��[�a��Z���;�T����+���gR˭,F9�w��x�~r˃Y�t�pB���l����~�:��p��/K���*�=G�vM���D�][L���r@tf��y��%I1R����`!�7���֗0o������T J�{v� dle '��kl\.O�k�E5[�t ��ۨ�ˉ��z��>(�>���ш�����������&�TT���*��Z[���d5??�$��t�p!��epӊ:�/�ֱCb���[���[ќ������r����Yf��g�~'��ss��*O  -�0�:+�<��Z��^�oOOr|���z��;0%�m�����|��T���ד�/���d`�`�|gyhUQ��AHD�
����{_X��<����|��M�i��Hz1@0'���I��~���-6����0(�:����ݲf�1��'`�x_�3�%#��D 3%����ˬaي�~�i���F@m%ɎC�;R���p^�Z�!@{g�)Lbq��)�J����c�R "�s�V��C��0Ϫ�m	b�/�@�@�@�Y��n@P5�.��cT� l'�>�4�k��'�W]�v�(���C�uT�j���h�ܱ���ぐ���S�����!�:W��������Ӡۻ�V	;��I?;����5��~q�J��"S��~󴰑�A����P�~E�����o4P| ��=��m�N�ΐ�q��=8�V�S��k��ؿ�зl���v*�j5n�#T�ǩBW��Řg�Vpp`m{���k�'��ME�}��.�|��|�w؍Ilu�s�䭏x�#o���:�]�_��'l,�
�M#cɺ�+mv��+2&FA�0���v�jh�@�14�]������U��"�ⅆ�0�q�<�oS����|��cg��B����	D���w�/�aW��������
�#��-�aZ��45����O88y?��8wnj@�q�؛�" �{V�{^�N���n�~�`�<���^N]kkk��N!���x����}��R��<<t�g�����jqlJJr���о�Z�x+2���n���eIq�
D�� E�c�3NM��fWW��;v|l� �Kߦ����u�(�nX˖�o���CJ�R�XY�2�N�o<|����Ttё 3�����@3��� �c�UH��|�MI�#Tc�-�f��#w������1�NV������I����s�Ͷ�U��ᇏ��Yy7(�M̩?��a�*�3�I��O~S-dz˨���J�)WK����
T��}�"�����A��s9jק��4�vIC@�ʁ�SZ\���L׮Q��H��j́����+4��g~˼�\�m�1�Vju50c���93��EP)'o''7>���J�2@Aن�[� JE��~�s�����ݫA�8�o9>:��=]�o�+��l?]��10� ��* P'�ù�Ӑ�W��ȍd���k�8~��P��Ic�����r��G���}[Z�b/��P
�� 9��;9i~^�N�Z�Ĉ��������>Hao����	��ۃ�Ji��Y2	=XW�wþV��q�L|)kS�L~�����9M���pWS�܃:���.��+� ��n��$�8���$�5�`������څ����Jok�
���'8g�w:T�?�Π˝�%j���4���N���F%�:a���ܬ���[^�n8|0O//��(����:(��5N2���3@h�H�;�*����:���a[��s0��Q�GÄ%OφF��g�J����? ����kV��K,��Y � l��	,�o���a816ZqѴ����v���)t�*
ID�hX��j�S�AK݃r���b���n�A���1�+����7@�4����yH�<X{���z���0�g����'rr�P�H������P���vv��߂ ��?_�Fz}��ȻH(3�'�d dñ1m����x��*���Y@�Ђfn�s��ppk�� Q�5�s�����KK�lɴ��׋*U��28S��D��%A��#���~�f�?~���w� ށ������!A��=T�
0�
��8��۞_�/�<7%:��IgC���6�Ɋ�'�x�2^T=ym>��r<::z۴�b���g�e���貇h�j�P����g��KH� ��RU�x��q� ~Z����M�c�
cۜ�+�υp�Gt���6>1V�j}��.}�]=a�I����Uo+���P���qPa :��1+&�~~���PJz��]]ݹ�O3ϑ���箇V��:�����w�! �K>��m^�JVRb1��llo7Yt���6��#�2X;>2���N�|���v�3�Q�[ݴ��Ő��k������H�B=�5eF{cZ�7f~'�b���Vg�^��[��)�/�{��[�'�m7^�[
�JP��<�Df���4j�lt��Ҿ�N�jg��D=�5��>���?��8�bX
X��_����C��b}������ �$k9����l�� W�B��j|_��)~��Q�����Y�ÄG��o�]��-Sa{���&�}X!־��KÕ�vxv�1�3�ԭCo�Q�[Q����Q�L���֏&TM��eٹr#�)0�~�~S����TV��2t��
�h�n�SqB���\TTJ� ���-Jj՜��.����-�C�4�7��D����"K�(����ר7n���X��-�OІm�����@�\\�A�����ly���� M��p��yoooh#U��)�lm(@�
.���t�
���
C�(��2��RΘ��Es�0H:׳��R����03\�]��Ó?>T����: ����3#ğHB�����G����-�k��TkkZ.㣐�AK�W1� ������oCű�'�9;�>&p���:70Ѽ�ϵ��l�u�B7t��I����ڟGx��p�J�:��%x����7��d|�	@�;ЫЎ@�I�K���EfV���I��;a����k�*����. ��������&�(���.w����*� n�pvgk��4G���wS�n��Uᜉ���241Q11�=�
�a,t��p�������&��H�AT�SκIL�]b�c��O2�s.��������H�4�{p��w_�������=?1997��' ��i?�4W���o��Z�%�H��#�?`�jy�<��+P����JaL
��[��*���ӵ��S��Nש���3_�?z��a'��������Rr}����tvwM��mhh�Ʉkk�������yM�1.�L��ӆ.��w�D���R�؍�+�m����%���'P ��6<C�끉}W���з�"��@SS3:]�w͖V�F ����!�XP?��j*��9�΍�c~L>�����m޺�3��ʻ��Z�9�o���_&�-�6+)+O��'���744uudffg8%l@����Q��ķ�6:���WD�\��ep�����6��P�V��R�3T߭��X���y����:Z���a)����5fL���0����8�&�^%̂��
m�9$>��cs?R{�s��V��ON;�����)��@��zQ���)����iv�Pi�2���c���ITT�9��옘�����������c�������l|z?Խ�qYRH���= 2�m�x:1 V�o�PC��$h����u���Z�� E�d�_������񝝽׸��'^�m`�:i��u���h~�t�C�L�?���։?��i�-�~�+�(�~E�JY1��VO���t)��/m׷�&��P`�ꉵ�@��_.�F��r� �.}ئ��o�%�@��@�yk�N:�k��]y�C��������k��0dB|k�6e&��~7sM�����N9 �|9�q�2��ep�ˤl�����w��b?�5.�S�*@\���_�hR3�T�����[L7?������r�pw��D|�����S6?1Qt?pCy���M��|�I��X�f*p3��o���'���1����.p������]��	�'u�ܱ�����3�Y_o��Hl��c9�Ċ��|q�A:��Ί��]���c�{�`rS�P�SMr��ȋ��,ǋ�Ϡ�H�V�!�U �omm������p����:A/���d�y���Q�F6o��`*���ｑ�(�X���dn���������9�}Z�,P`Q��
�� �;��7F�������B<ζ��SRRn�(�������c��%;���ڀ��Vș��Y���6�p��oRp�>Z�@D/���a�kV�frV�;w8ZעWƠ���<f��y��cb�=6��W}Q�M?,8�h�HB�$u:6��3��_x�*���ԤT�6��9��A0���]*�`�T��h�����@�3�r�@�ж(\�f�̪]�!N�bv?�I4���5_���=����v�T�.-��s��1����9?T:
�Wl���5D��k�^Cc#�U���Ufqfff=��fM?�Rg���#�~��lvՎ��՟���t+/��:��G|�o�[���!b'k9}�=�eU=c��j��Jq�c�X������OLOg
552�1�����=$*���K�$���Q�K���)޴�՘/I��sT/:UNUxz$�?�377E�B7��VsTVX��l�jG�������g���sq����[[Em3�sB����:&��7���Q�9�C�@C�p�j9:>V�C����}��h�X`Qf��c����<��Q������ă���\'�4&���������x���ٽ�1��h6�w�ޔ��g~�����߳VU���7w
E\�5اlnn�O��h���@Y�C�Tyi�F<��}�ZY999�l�G���O"��%�+�F�摥cG���T��J~��YBozf<��Ϙ�y���3�qkL��烦��خ������2l��oSxW�f��������LYV����V�%C{���s��s-E{���A+햷�8��s���S�U��3��������+����%�
�''g�R���үb�%���:�f���W#��[NMƃi��z^�8�M�CM����S}��FyAΞ�9�@�|ms`9�ҿ�-8V�^t���Zƽ��Z�K�΀�9Ѐ]9�I���'}+�g֙ŀ���+�f��|_q���*ooG�Z	�..."��\�d��%�3�{�z\-���yҜIݰ��6��$��g�G]���iT� >�n��5����� �yG�I�߿�<�Q��q��z~

=����i�j����7����Zo 9��L��n�_�o?�ӥ
e�Q�?�z0I�G�/��������eGkk+�i�Q�ؒ�їC�[�}K{�4 ,��/�ЦU.H��^gr�{���c�����=�M�T9M�3�ͤf���t����M�7\��j�}5�����a�䰵�uYU�V��
=M�T^~b*�b�6z���/W�gA�y�;��`�'��4z���i��Fa�D����z����˹
��1C������,-����Jf�(��"- )7Vc�����[;�g�g����:�lub!ߣV$ظ�0�z�{��-��&�9'���ΒQ24J�yZt�>��12���;cE���2F�V� @n��Y=	�|($TVS�yu��ЕE�[��ϙ򦁥�:(S[[[�_H�ek[��@��\(&���[��@�Kl凜]wou��!��i�<��w��\vB6B�xn@'��HB����^������b���aV�Uz{�C(�\9���KU��
��+���u��j�|0+�.q/���B�k9�����:݉�!��ϼ��Fr���@���wa���u�a�m~vw���
:ϵc���F<{_P CAA��� �z�8�)h`J�uZ����p2@���u�+ukM[��<�6V���UX��=�J�?�<�)�M�ϟ��@�&����r|���Q�K>�-�i\�B.�"����$�=�	�^~��Dl���,^,�Ie���}��f�|�V\�	�c0��گi���ܦϋ��KoԸ�;�~�Gi^��~�|��Xс;�8 ���Q��� I�Ф9�^>֘���>h��P��ܝ�����F��U�p4��cL���Qٯ_�b�KU�7(����By�:�T2�s�p蛜�w�?����Er=�)3@oAiv�w��D�c@�{n����������x0j�eH�4@��ԋ�ܜYx��묟�ƫ�R�F=c��;D���r	��t6���j-;�q����oҢ����4ϣ�a��U�۹�cS�`Ri�ݗ���� �)|�R��~-W�n�5����(��峺�v���s�%k�"#cc��k\B�l��s.�l�c�8Y��u*�P��.~69�[�U�~S����9�V�d)iiPf ��;*��l�A�//%��-�	��ß���T6�A5K%v���6P����A���ZU焻R.���`�w��^��1��!%�c:9��C�	���CE�T\��rA��ކ�5%�Q2�������vߣ8�?X�`t��*��~���dT|��s���
�CpnJ�bod����z�D���4��$BMB�
�O��S�UM��ߺ��Dn��p�z���籢~pj���K^�NqT��z�	)ݲ�����.z�Ey�辜4˕�k�x�5a����5zU1�$�=<t������XR�L ����̲6ϊ����蟼?G&�WK@IFūA���b�&��F��*��\�m~��~��xQ��-w�o ����ٿ��V���v}Lļ~�w��v;kț����o�:Ď��e�5��@B�7"Q/�h�J3�["�Y��M.��_L�ݮ*u��@6{hp��Td��_�D�Ȕ�ۇ=�������⟘ӟ�*�\"l���J4��a>�ք��mU��G[HaM�j	*�ѽ��_�����34�̪�ǰY��Vm]gb�tk�6� 5��?�_�]�'��^���d-����T���L1wO��Re�.�T�p�K��Wm�;���~��GNp�f2I�����v�t����ᗁ�v���~u������ÒH�ƃ'DE�ָ�%�P]�j��0L�1��~��D7�J�4�y}^rU�wf�}跲�c������˷���z1��\Ͱ=��	�A���BϫV�]F���e�}��m2���-���kcb�V�%���0��3�(�m�4������i��#yM�Pz�������԰0����kվ�*=�j�P���sv98�#�<��O)mW�w]v�G��5��=�\�7�%����<;ޙ�@�4x���C�c��� ڵJ�{KC3����38�B5�rļ9�v�Mf���I�f@Z��k����*��8*��d������1��r*5��0tJ"pbzU�8##��㳛�ț}|��e�w>���@y�?]��/J��Vx~������[[�|�〭A�^��`-/�l�}?�>�@����4��J�߉a�7�#W�ԃ� d�*�V���P�by�~ˈ��~��[%����ܐ�7�z�aA;݌�Ig�W��j��6�ʰ�Ȍf���Ub�gvB)��,]��-h{{n^�!m�ʔ���6����������+��&�K��m��J���K���3��_� �֐���qj�l��9�߈�J��S�����Br��V\����@����i�o	R�����1�{h@�C���������V���gn�E��ۋ�r��_�SǾҸ8���,\�A�}a�W�ȴ����u$йPa49��;�w�)P[�j�4V�;��=�vC�83�d�X$�t��4�m� ���''�

*���JUq�����7�;�����E���n(��n+&I�#0۩~�����>G?�VH�qO����>�
1�?�ׁ�K�R�iv<|"��4�ka"�8��z1&6Q�(EI� K\h(�
�O�GԒ�V�t���K�wrw��z�TIݶ7�ᨋJ��O��Nl�yLOm���w@�x|b��r p�&Wb��4A��0���q�ʕ6�2X�����t���@jL@Hkjj����V3����ѱ�O&�.�(�Ǯ"f��t%"�ľӊZ	�?'�b=�3����+�3G!ۼ�ڭ�Ɏ�S�c���1m�Pxm��cgg�5Lw}%~
���}f��Ѧ�;����iU[�Y���v����?A`p����C��;8L��U0��ƮC�rzz魭-xU�_��}9�o� ����2u �B���h�k�x�����`�D�//�5G�{���bR�XG�)��i��p�f� ��F�����*w2_��ZUg�8�Z��� owv�~]s�����G�EZP
�����&D_	���϶^��R�;���?A��7�|_��Q��<����Q���W�cp˻}��w�Ӛ���@R\#������ ��C��(��zc�||v�z��C��R���7�T��z�1_C��^����7wϯe��3N���[��w5Zι��Ҋ�A6���(��<����{�H
�&�7��:��O�/XR��� ���ŋ��A��&Y��?�҂<�7ea�>jr�i.�� T.b���O��q���y���4#$$,���pa� ������<)��ќ�o�m˞�6d�ui����R�xM�~�@+���%��"���t�>�V�/�lŗ���Lڶ���n���]�R�y�g;kj;n:�E�c�Ꮵ;O�Sé*��ٕ�|��k��t2n�sH��Y�W�tݔCf����.ccTž8�#%
���u����x�k�μ���Ey�O�_w��կ�Pl��;J"x���[(��6ǳ���?�r7���'g����ߘ��m�93���L�-;�؆�ӧOߨ�zušZ���)_��bzܝ�r("	c�-�#�W���sg{��^9�Zv��-RRRBF5��XkC#�����j9�����F�P*1[*���bS_��0�ޠ@�m����L��fr ljjj��g��uj��&�������c��lpn������_Q܃g��Ni�d�T���j}֓sC� ������k��S=O{��"O��P�msZ-�H;��n�1o�)o�I�53^ll,C�
#9>���e&�RY�gƲ��{7%ɲ�PK:��t�J)���uT+�h�OM���AC��U�~��m�������kW��֖_@ ��/��#�O�/E�\E���:&H(��\��>I,��UQ���Y��Ls(�=��J�R�������i�\�M�Y�~��e���A��~�t�6�!%�L鎂��vz��g�m�u��mCرv��T�`��2m��`�5۾�+��1P0�1��� ~O�f�C�+�*�H����V�n5+"�a�e��F�+z��]�ӹ0�X�Q˾�@`wA��n�Tc�͉�!��-�ҕz� aI�\O�������Q��ks�\$�T����b�<=��ʺ���~r�/Mŝ�bV̉��n�ڢ�ĳ��Ӷ�y�ć���?-�Ҿ���W�.p'|�{�;xCt"�$L��r�<ԋ�~��\��N�~��hy]�g��A}���o�����a�s�3�n%2b4x���7Zg�665�ttZ���O�#}���(���/��R�f�!h�~t[^g=B��d�'��_ؾ�L*�}>Y����0~�┑9���X�YE*�KO���-�_��UFK���������pS�"����204�98��Y1i��q�vh��Ko2%�<��=�An=�� 1�˖�i��f���0l"C��]F��:�g���9�К�>{�7�$~�	cA!i�e�<iT�i0�p�!�I�pO�Q��x%�'�2k���զ��$�R�YxVz�����
BV2O^��PS��Y4Mp�T��7�q�{�,�od��fTIiT9�$�-م�A�v�mUeˋ,��^��`ꏞ�����.{�`NF%������y���z��o�1]��#��"����9IhB�»S�S
�I>�%�u��A+���9��f���2O^��˻ h0��V�nX<�D���o�
�Ka^�ċ1����>I�{WX)�ݬ=�]���^z��O�w��}���q��!o�fƵ���b�"�τ!��ymy�-���� >�*�W�X9r��e�����\E�i�\-)�_|����>������=�5����ig2�z/���:�1��+O~la57E{�JT�]�sX�/ ������:�>W�vW����Mے��
�`V�<'.��������Kw�����m��&��xF��2��J�zJ���]N���N-@��0�����|?���#ؗ.ELp��;O5e5�[�Z.���".:�I�
��:<=�{G��:��p7#��`>[צ�X�_h<��˲k;��RG�x&.pA�]�U䎽�Ӫ�������c_'����M뼊dV�s(ܼ���(��f�a�>�Jmd�Ã�!}��m&�t�	�ӷO���e��'�uu'���,��������f�b�_T]'�A���@��l���I]N��x�y�'���
gN�u�����wI[^^�o杻���ΐ��v�>��j�VY㘭���=��c�Yu��nAU��C��.Ů-��[�n���K3��Z���0d���E���M�>�/��T�ݐ+�#���DKg=)��ʱ���00���ĥ!��km��8�m��=�B���^h��=�}������)�ﺦ��e>��M�T�4��x�H�_X���#�=1|����?yZ���H˂9ʲ��.*b���z�H[[[��
��0A����0Ѹ���>�ّFˢM�u�n�F6�����w
��,F� q�ɻӁ�C~���13c�,b[!{�|
���~�]���Җ������)ACG�zZ������o���b�Aھ�uӲ��҅��=QQ�M\���G2_�hlo#7|%v�]Ò'�{f���Zt�I��L�����p/DW�V��E٠���ǟi,[`�;��<�i�#ɚÝtg�����i��b�O'��6C�����Vr�ӣj�-�H����R��Y[c� ��:������J���������Ғ܏�_S�Y/ϖn����V�)fWZkpg�������ݶŶ���  ����<q	}_s����
�tɨV���)J�'��|�{�9Ue�(	.���8G�d �)f�?��� هl�v����{r�`�Y쮖K�x!��H���Q<p����%���ka��)������;-��C��M�^t�|�� ��G3��aJ�&��b��H��j����p���3nv�7���$��г}�l�5or(��6��_`X"�B=ww�ellL}�v��23���Y����c��O+�i�@z^�}�ЫĿE����-ڀ?=8/i��nɼ5�tww�g�.�$t���cCKC�� P�"�R�9�Q�G[��I�^�z�Sqzyq�H�ENqߔ��(�Θ�Z�V*����(�\�ş$U��-!k�����ڑ�d����7�.*����X)��+�4̜�j/Q�
� ��ҏ�Ҳ$?�ׇ�0;5��M�ԛ�`��'���V�R�-љGeT�+[p{BlU}Rчe��m��n|�H^��J��O}S^�(��O�\vZ�����I��r#�֣p��i�6��ٿ�C��?qJ7)�{X���y��}�����*�=˕��n�w��H�84ivA��x_�d�=�rH�g�4���j�!4iqþ|�/$$t4��Ԧw�I�݂w�6��D=N�Wf�?9q�����x�/��5��2~ϓ"VE��󇎎j&Z���������j
�6ۻ���.q.LFd�2a��Z|���_��
p,�Q�Rt{�Z��w���{r<cn̸~&gܼ�[�Ўݏ���S۶w��%?z�	J��[_�q�_��d�h[c\T�y�q�`a�T���)
��!�x81e����B�|>��an��#�-�#�z���pU�ez=Fا_�m�ުZCwAw���r|�Iد yȑ6[I|��c�>ߎ��}G���n�3j��zOOE�J�Y���J�U=/�4���A��|�b����>%=n�������RVVnv[��2����d�.Ցʒk1Y�R���3�#��(�^z	1x���,a�J��x7v@v���$�.�2��}��M ؅��
EZ@sI�O�1nZ{o'�ƿZu�n�E��@B/��mX4�E���X���c���ؤ�� yY΀#i�,'����4��|�$�Ik��1b2BsW�HR�
4�5��Y��a����٦�5�"	�}/�H>fA?�H^�\��l;tz���?�6�u8�������p�gMz̚ԣ|�#��v�-���{b������������~p4��yUj�{�^��x��;9;���9�
�H3����ē������Y ���O��>y��	:R�����tz��YͰR5��K__�
k�ͨ��E���~�V�]�	ь_p���,�LT�@�t�m�B�*n�I��0���-Mw�88��q���Q�V���Q�^7���<��Jw��v�������P�?}ɋ�in�e� Ģ�"�05�U+�۟�����=�� �FC[h�MMM�P_�%��=�H�t�P����`t=6km#y9�@��o
צf��T4�KWQ]��ӐU-� ����b%j��B¹��[�Ehq�bTX1���� t���sIO�kҝ�.��� Q�OJ*|�	/N��v��M#���bE@P��j���i�Ċ��{�z��M-6J���Ñ�8���F+3���i9�ݺBL���������M%�o��%`��wc�}6:n�����e�Fm�`G��0�e��ý=�_�>%����Ҟy�R�~����$�Y���ݾ�5hn��m?���q<ck?[����������9
0�e���cwZ�p������X��1/]�>�$CL�8���w�4��K���3�ݕ����S���2�����#Tsgc;F�N�-MP*=�R���S�hr�ѫ?B���ho�5h���Y�1ߵ�ӥE�'Ѝ�h}�[?e���#�@K<�H��S�.����g��~�w�l�4H�[	Dd����ѝ�x�qy�JF	������4���w�f��o"��4��J��v-�5w|��mN� �� ������{Z8z�̽�a�������E����R� }��=�qooO���N܍��»��l��K	RDh r���Ax����-.jݩu��_�Z�fIF��w\�u�+9ő�4�wo��D�����T��]K����F�+־���4r$���T����L�f�z��~�bbܦ�] ����p���qC�ZbACMU3�(��Qc������F�%�i�i��~�◔�`���ˋ�0ͳ����Y������;��A{��kǙ�;˧��`����E)�jA�J���,wq�j�k��t7p�3��)RA���V���'E���6	�g;]	�KPa#�	������*+m��#R͝�F��U.HU�2a���F ��47�G߈ ���;y���Vm�woe�m��4ޏFS0"���~�ES�<¶jSS�k��Ѯ«��)������9(2���$��`i��}'_q���M����"wp���ʟ���hoTX�����|��J_������l[���~������ ��M�Շ��P�|���B�C?:�ٟ��V��/9eq>.�-���ͤ@F�+��wz�:�P�����9�y.�L�S�]>��0u/:�o���R��� �p&̞��.�r͕�a��l���u�)<ok�G�Q|��]ϙTzQ8�w�=_D�A����.c�呋�P����a��t��y�Yr�L�q��L���/_nX>����3���L�0ē��4��*K/��:55F�� ����m�Y3�.��&�;&D�|��������s��',ͱ�5!���j������������^]~c?�/j=Ԫ����^o0uR�Ļq��5?��J3�p���\���~Xo�l���M�R��Dl�GX��#��q�܉�g)��pzG

5
�jy�v��a�3
�5r$���i���vO���H��b�JF�e�>�����X��~��ٶ�}K��4��c�9���CԔ����wQ�)@#66� �<�MJJҘh�Im6G8>��Z�Am|{�*1��6+9ײ���F�^��ZMK�u 
����=�S����~�;	]�G���﯑��Aሔ.��*vr� ���@���<a��0�(����~>?w�k��'%�?*Xͪ>}��gAp��޷��#8n�h��z�$�/�5��������S��۲�L�#dI���.e�p{^Ua)���y��#��4;x���㛃>�]�m�?��@���*����O�11�7A��k٨�&���YZZ���ׯ�@����;���5w���5��VcdO���Nf=o�4������p��7�/��7�m��Ode��UF�(a�h�=�2a�~�<p[���r�|�*�������.�]O�t��Ԯ#�q��rȤ�0��0�Q��/O�ʋL䬣XP�/`|�J�g1�����90�7G;!P N�����#%N7�-�{P&_c�\��p�|β��1�e�Bg_K�k@*@S��k5k�bJT����"+�����-xp�rW0K�q�� �'E���Z����ڑ��S��࿋�3����A
0/�gN6
�s�~�ʇ� �T�+e��yX�=:���&���C{+9)a�&ME��A�p� ��@,�����#a�	~����^"�����0�b]��$5�t�I�q^�����ˑ_�4,�@��q&�{L�����1{yNp�"-���R,�4��^e�ؕ��("�u8pv��0E����ɗ@v�n���y��f?�$W��7x��-��(n6�z�ߴ�ϭ�܄!�[����l�C�ڒ��[^�Y��G<9�:g 3jk�cT��d%��X3�m��M]Pߺ/���d�����9b^���[QU���w��4��	��r�X|B؛�L�]*4A��.�)��W��=U+o#nǸ�?z�)��4�������S�p�ga�z� �ג�%�:Q~o �j���s �,�f�"D�4����p��S�a��dI�l���N���6�~4v��+i���l�ͱ�d;:��jB��0�P��h�6�D�ڌ�ӱ��z7Ě`#�y�j:;��c;���9EU/	-	K��k��91��9u� Q�0�q7@�	E��?&`�ilaD�%��2����[��H�)g�铙��Kǽ[��t)C�ϗ��S�c�d�����ƞ\aw��*����K�s�.����]�a�����	�	����9�u1=-��O �H��2v�_���F#S�	c�[��%T."#�2�v�{:߿��syq�;���9	�[EU���eo���,�����\X�I4��x_�K�Ձ���	�my�Y5B��XY��x�qw6?8�C8�=uF �����j���|_C���_a��D�S�Σ���E�7�r�|��rn�㜻�?a�g�)��E�]��2NAUw[����������3�WӦ���W�檛}�G�mr��7���p��2��mghy5E[	� 5%�!"��}��]�bͫ�.<�}S�5�����-���M:ڿ!�q14�&��
�"�S'UG�.��zwl�n��a�<$d!?#����Y����`z�5����E�����O�j������)���=|S�O{��v��Q������0��u\`�a���/1ȓ�F�y��J����O�rް:E���&�{*�bee���A��窷�B=����6��� ��-����0˥n�-�������Ĩ��KMF?8�C!��S�^�~�Ǒ	L�����둙5�l�l��(��[�M?3Og���[�l��~�wr/F?���D��\M�\,�i�<yZ�=�- �m]�{���p5L嗐:ޔ�ì��88ǘ�ࢧ�*1�%2$��夁S���kl%K:rjqZ�#=�[3`��_VD���ԡ7A|u�����#��Qү�o�]!?YO=��LH���R�7\�3���s��,I��ȕ	N����u���Fo'^��:'����miȎY�?�A�Hݜ
E:���/����q8y��K��.�iW�8C��5�������Wܼ������W��_�x�vǹ���.��ȟ
ʊ�7�F�/s�����\�A�_��V�/�8)c�c�%<��}��@s�S�_����?�aA�T��w��j�X�����9o��>���h3�r|O�Ry󟼳݅��j��x��KF�*�1���n�I,ݿC"�w�jM��KL��1k裠j�%A��| Ճpo���dbbz?a��{��d
'Mu�:�v=-����y�Up���Be���_ǡ��Q�X;gPԐq��9}�t���N1��qȣg@��#�� �E������Zn��=4L�G�z��9z�R;U/"��"=���	��(wFg� ��X�mX|_�6�{��B} #��y���������G�0�cX��p/���Oռ�iܩP�oݥT$����� X�!+�+����qj�4����������1���8�jÚ0�,_"�R���K������^�b�Y'u�6g���d�
+������p��}�Ju�� 'g��+}q����57w�9��(��)!�}/gE��,@�Wa�M��9�(�h����
����mA��PB��.IA:EJ��;	�Nii�.�����f����{ν߿��yD�k���;��c���n�P�V���j|�f�Q�3o��[��n�5Q��)���R��fM.|��=`H��nŘ�t"���4 ��*�|�G��Ls,�>�݋[�7��GQ���*��*�tO�Տ
����|D���K��9/��/�?�`;Ra�'.�P�ޗ�D���iJ�p}������c�_J���-��rw-���sn�T*��z|�[��}9cj����OP�ж繋�Uo�:�8�A��y�İP_)�,"	I]3��4d+�����nA�D�G��X�`tr�����_f��~ڔIs����BY(u�t,�%��Z��m*-�-)�Z~|~ך�H9������U��9�,E>��r8K)>�l��H��Gt�=�L(?!&)�����+P9Ej��,�����tZwF���^��B����A|��P�r��G�����Nd�n}��B�l%֒c߬�;鈙jqFҎ_FOA�E~��cR��x*�~�2b�nt��@�	�N��ӻ���k���X�
zlu�goh�V�A��I����{|e������Ajʾ�D�A�~D3���+M�E�3S����AO���m%�Zƹ����y�U$���ʋ���/7^�"��5 \�!:�*v�C� # �����;�*{V�;��%z�<�i����{�F��0&����E��'KQ"�����r'��1�'^����T���!"�6F����bxg��h�ɿ<Q�9��:�����J��%��X���̋�̋
ĩx���m|i\�G9�+9����ɪ�b�5߬�����OD@_��YJ�1�7��!�W?L�Nի:k	�g"�S�Ey,X7�֝�-�Z�g��;��1)+18��QP�q�^�+��j�\���w��P�O��5�����^��!m;�/,,��N�Y.#]:+'�<�g���I��7eQ�o���������,�0���R��l��`���Y*�F��e���󓮷��Ϲ�;o����p	m�u΍�8�#h�v&8)�����rB��Q��dkR��Sw�D�b������|�jM�Oj:!+�{F�����]��uv�f�_���ʨ��$�`S{d������#�v��X?LF�2�y^�z]�	(����ῂ�-NN$3�S]=}N%V���x� r�h��sN�4p3?h|��P��0恡����!�H�!��K���$�i
�ܝ��]����	�WfL��L�2]�9��=%�R�Z0>)#�R�S��䈼�{П��Bo]%u�Ͱ����8���wS�
��r���(���e$���p'�4oBV�/�X�6̼����{�>���`����6�3��M.���y_Jo�?-TB�1`F}����w�=~�|\q�9�&��B�B�HK�y����w��,>�Ǐ���irˏ{�}��[I���h�ŗ��~P�ex��"�]�����{|}�z]h��55E�o-Z�o�[����C�nP ʫ���Mȣ?iqpz��z��f���hJ�a*r}ٝ��@o���W����r�6m����9
+��)�$c+Ϡٟ�4�5�Va}Bq"��E$��Ե�&jf`�u�;���6ǌ#�SE��v��������l���]J�ٓ���hs^�]ى�Vz��Jd�N:�#�Z�GR�@�Z7�q�}K���������-U�bQz��$>���yK`\=�|w!��?��[/�(������E��S-��H����q���M�.�[Jl��yq�g�m^�xw��rr�l�B)�Q���鞢�ڬY���7?��H}c�U�.�n7ts�%�{з�[���J����b������i~��=�?�ٍ���'�"h�9�����m_�?o�񛴚�tR5�ҼY�i'Y�T��[-a�G�}�{�CN4�y�	��^���0���CAz�l�з[�q�����M�j�0�\䲋�-r1�܁3I�᧔�f�ժg����Ab����x�OH!8~��|�B���Rj]&\>w8ؠ�g��t��L��ֲ�6-����ѦxiQ��o��˺oM��Y#Qb7H�f��y����Ӕ~�k`���&��F�^6���:����#�C� ��- �\T��u��66e�Jq_���|�cT~g_0��}>L�e�*sX�m-4.k%�!����V�f7�l}���	f�ͨqy�����������R�g-�L���d_���˖���|R ��zw#� �y��Qv��]/߅�q�M*'�S����W�d���F�*��_�А.�ݘ��}aƻ6n;}H�����1∯A:@Aam�<́�&�{;tXd�%��s�����{�ƹa���9��X�4�cr�+��e�~�@Zc��ZL�鼝P����}q��;%*5��\:��'�4��*����J�����mٹ�� �t�i=t�_B��*����L����$�����O]q���! !�*$��{�qu�H��&B�sU���|�����V�1���*�l�I܏���_�����zC���S9x��I�����3`�Jy ��V�~ŜL\x���껵�sQF�>���
�P� ��["��i�H@�:@��� ���ok�M�[cߺ	F^(����5��Y�?��D�mlI_�joOw|dܭ��yY��A�[9�nC~�=��R�,��b�rcIf��##8999o4���n�^��o��~��-r3��B�|r;LZ�ݾ�8x[� #��1�#Q���t�*e�_�7��D��Vm9ݽY�'�C�g��+�wǟ�`W��0�o�NTy��s�7jp��`ﭷ��ك�򞅄�9]���b���f�����"[��y�f��ܭ�&{<�J�� ��Z�>�+3�,<!	���ߐL�<=͗?��� b����kk�%�ߩY�(�[���6(��^z��Ͽ<#�G����|�Ԝc�?�������Q���f�?{�6L���ð��
�G�D>��+�Lh�n��ў����֜�s���<�����������0�%>g��V��g�FFjot�`޿�����bB#ꓺ��1y��v1���)?�7x�yx�L�:���������#MM͟�~��L��"�jHd��]P���32Ύbb��>��Dj��֜A$�[j���>|��ya���]�
WW�.���O�s�|��i���QZ���L%�_���\'�*1�7*F�vu�͊:��o���`X�+]#>)�ml���s��X�ak�
��Uצ��T��_g��Fc8-_R����8ߘ3<Os���0�K��_�
6��4���]~+]�hh	oO=���9��G�}�A�n��d5$fܲ�����s��e~���I��-�a�^L��ubb�>�@�/����.$��پ1z����^�����0�!���'��\�x�n�h��x�u��O�ש~m�Zu��gл����&bA/�%�n���ޛn�u������x�� �K#�{W��~��9�� ��)j^��P��^fz�Q� �t`����b�d�$��]�����Ꝁ(��[cI=�>�>�`È���-�\�5�j�u�&�h�߫�y�.�R�������1��0�O~�?�vUa�ɢ�}�l����П|��5$�Y���ǩ���Z����a���l7�Wmyll�1��u���Ʉl&8
/J�B
��K�Z�N
���ОM1�C��8=�N���*�*e@1'66����L~����'����v�d��J��<�9�)�OR�F.�/$��&�2>CF��ZU��;���W�]GE1,��ג�����Vc@qJՍ�i�H��|*�����;ґ�F-6��27���$	�Z_<���r8o�=���L|����)|�O��F���f�ל9��Ny6[^^�ފ%�5)?�իW- ]c��ic�]u�^}�j��9�+�|�	~�E�_A��o�,)�M������'$�N�|9e���C
'�Ϙ:6�V���ԏ3�~Nj�z�Pj>2�'�����5�ϳk��WR�}3��++��J oD�;J���A�+�$�S����
ȗ�ΆJ��û��̓�>Zك[Q�)F�o�ghk{�fl�_�␑��A1��?��)�sl�� nˇD%��Rk��ʒ�͚=���%;�O�.7�D�\Z���A��Cg��q�Z�����̎;��^�_v���~5��n?�����tHuq�s-����2��bTxVkͯ�fه���5���4���ȷ��GR�(�+;�ʕ��(D��1J=��ǲ�g�U�9�.Pl���?$*/�ǆN�~Wk��fY�>��.:����^��F�_Ϭ��Y]�85� W���η�8 \I�,'�Ő#_��j��r��C��-�}����a�=����/F~��Sf�$�~/�y�����; %R��D�qӝ�k�����U��PO�Lb��p�{�wB�J��. v�φ����て�=흃�w���������J?g�н����Sa�a������ѿ,&#V�����0���f, '~}�`�8�)/�8 jV��.>���vz@:���[�{���㷭~�[ʑ
C��'@�P	�?�K?�~Hw}V��k�h�c��zy��u+����c��ϻ��U
TUhq����,��F��oo����$;|�����l����/ip�E��qh�Iݴ|�լP�����z��r����C>
"6iQ���g�q�>G{�w}��u���E����	ԣ1$4t��.ue�;P�!lU�� �F�t�<�u^�FݟU�ޕ~��\��YJϲ�M�_��;} �:d!�k�X�O���:�(
ɓ��A�<(Yf��x�/��Y���ͽ��_���P�����u쫻~\���	��͗GVל�����m-���n���A��������jam9��L�a瘐'���H���5+�{����8&ݎ��@��ϝ��K&��r����[��E��OŰ;�=\��X3���?v�M.��������0�~�հ+4y��Ed�f�'Q]o,-�߾s4 @���
�Yz�1a�� زR�-�XVV���;`�3o )�&�/�Է��㣥:�=ҧ�/O|�O�ؾ��Ea���b>������E��_��ϋ$<A�c���he�F�w�nB��98
�� cvW�%�'�������TH]�|[�\�g�.
:�r�����Df�+��8�<���Ӌ{mn�T�E�{�h��� ������<��x��)诖�ުW�M�� }(��q�?3Z��}|BpWp`����Se��fBwۘ�VU�K		��?��<	��SA�v0�N}���nZ��h���C/����[:�� &o�|�*y�o|���������v��k��_�&���P�w�P�}O�A��@?�,=��V�L��o��m���
-��ܽ��ݰ������`�N�ZX|��s!g{���Н����9%���_�KK�iAؕt%����n���tJ��9I�9%�h%����j� ,�+���f>��ф�����@��L� d��.+$��<3�4A>/�ߺ��m;���QY�FT�ڶn?�Ǘ�$����DD�?s�������KS��/�۽����Ĝ9��Ey���%���>C <,,,��#��O���8��'�ֿ�8��"���� �HuF���>�Ըu�Faq�c�r}�L�n��A�kk9�F�y+����T�ҩ��gAF�m�`C�$��Z�}�{�e{y� �X�`?�DUiSShQ�\����4ϳg�4xxx�/(��� ��o�߷��T���r�IZ7n�6Z�-E��Q_#�[m����]����t�M_όg2d�GV5�s���ǌ��4�+Փ�v_J������������洈�����:�N��d�� ���	߼���,!��ܶ���B��h9�Pp��ÿ�{�N�5�j�-�?m��\ku ��Ѩѳ�S��v6���fG��l?��M�ɻ��ܚ�U������ 
�dg��1���U�������-7���U�Tj�M�u�[���brb2�'l}��4���X�z0�����8�U�i*
�~n5e�L��NQQ
7��z��@�؂ss��7
뛛�e֩��J�'-�)��󥷶����o	�>ʮ
TN�9ٕ�v`�sKQI��n�<k���՗���oa�3��	yƅ��Yx��Pi�t����S�j�;m�#�Ù�����.�_���hj$�ߓ�����}��2>!Q4+���s)�#-����P}��OB����߀m���F�to�ȕ��)i<J�㩬�;���C�������/��mm����]����������qX��dd%K����?�����PTW'w�D��4?�V`��CS3��Ǆ����~U�|/<�c��������O�C����WQS3�np��G�k�4��"Џ�m�"3��~��
oߔl%���9(���f
N�:X�'�:ɼ�m�)#^�4y���G�%`�:9�AEE]��^�O�%l��IIIQ��4{ Z�{=��?<x'[DE���ӿ��$#*ټ�֯N����0P�]���c�����[Ӎ�/� {�ʃ��\t�grnd�r�p�y�U]�o�-0g��2F��R�ƠWg�ƿ�"<�~�ܜ�Jf2a�	U(�
ϡ�)�����PM�u�]xś2���DEQ�I��|��pܤ,���F]�x�]S��t`i�OI�x�����)�ŭi�&czP�����"y,wE����q2�є���#yʶ�Z��5��tt��ө��V9Q�׸O9��jsE��%�ћ����>o~?Ӆ�6������7_�iV�+��޾�N�R���.7p��Y9��~���� 	���ò�e����'�t��̀n�B@�~j!�4�V���@ �?%��Tڰ��%TǪ��c��PV��roB"��%�~�k�vQ�3���&�(���r�9�f�Ak��/G�N$��y={��|�w�;"�38������d�C�{ֲt��d�"�^2u-��55�D��n��L�K�s�ԁ[�����(=���[���hQ��F��ߤ� !qty�sN�+ǯ���|�<�R��ow��m-ҾB�A>�^�,۶�P�Ϯ��p�l���)tT����~���P�Mm���D!/O;v..��4�XFĚ�ģ��=����8Y8>UD���}��k.�+h^���e�9�Ɉ��]+�<i��:�%P�X3��F�"g�P������r*��6�2GX����fҤ%p<�����U�Mî����{���Q�ǋ�C�_I^���*�����!�V�i��h���kn����ds�d����,X�h���_���I��z�óU�`�\��X�9�mS� �����T;*�A����*2ى7J���ZT����@ l����/ϏW���ע%�N�`]�E��hh��Pě�������-Gd���^?�j��~v
>�6yN���Z�KRN�i7h�T����]tvvF/)Stx�W^�u�v��4���o���
u���F؟e;��{����B� WLMMm9w�.���J�̛�U44X,�?uHj�����o� �W�V��`vS�oh��Xt*Z����^�xdU���a�1;��ym�+Jy��T$ZK)��P�9`��[p�J=M�$�Ϻ�}>Ł����Y{����3=%��Ca�@y�������Z��,���MoOՏNM�T�j3�-��$!~�ў�j��hOF�d�c�<Y:��8h��p��6���m�&��B4��G�{��6t5��1:&��5���gN��w�c���k	d~u@��p��Ҷ~
Ec�]���.�99QQQ����f��!�U�/_f��d2�"[o�x p%����@��F�s*�L�#�'����4!�p�C�yu��m��e��$��n����wX�I��ן��vAi��,MEZ�C>b�Ps$38�(޳s���1̎����
��:�I��x>�b�Jy#�yϵG�h���b�P.H�u.���p�����T�[�⺍�j��Gͩ�KG���N��^��Ed�	���k�����Fv�%�Y���Ծ9 �LMT��o�6@ܤ�ك.��W,��0+v���Q~N���1��/�&F{]�o����p��&����G��s�	�'���:6�ݎ�<���ۡ��#�
PJ��$4:���A�p���z~Pf�)��c���f#��&��/��>)�`�=�|���)��r����u{��PY�j6V���1N�Bg����|��]���ڭ
�������I�z��ı�8�ס����D���ͼ˞�z��������^FO�I��pbB
Vt=��&���H�_ϋ���􈃟���̵`A�HSSS.	k����<���9I���==�	C�R�{���DYR�~��3����-���xH���Ϗ��@Hٝ��V��(-�N�O1�<�$.��&�sMM>3K���z��X����.f�+�b��N��<6�o�ҝ�Bw^@7�A�i�e�U�L�������{���+tbד�����S��4uX��C�A�\n�AUTW2̢||dr2�Œ���FL�N����w�J�c�<�",�����Q��o	��C~f��g�xA+�Z�3I�lb�Ka̰:5�1���8qC%X��絍���cR�ۄd�?)v�n,��,^��,i9���o"Oe4K�Y�a�QTEE0��6 ""RQV#�����Dz�g��$�|UUUt?�Opʀʟ�ϾQ��%�P�^z'm�i��^�zt���G��i׿�7_Psf-.~�l}��4��2�G�g{�Kc���h���/�k+� ~;FE��S��ϡ鵍�њ])�nk�Z�3�?�a/��� ?��r��A�+ �!�556��+'g��T��-~���s:)++�����%�;���1�]�#�u�zrkd���Z���_&����Y"zAɓ��0q�m��E�v���P9z���t����z~�3��Sn�v�E��`��t?�R�S�9�\�PK&�%%��I������$���=��嘘<J�Q(�z�$�<k��rHN�h����
�������*��i�-�%�c7�^^ƀ�ë��� U���hm/peI=��
''�Tn���9y'�,�a&�0�AU=�b�����zw���|���\�t��7�Z���"Ǹ�^d��u>���?���p��9󃠤�ht}���ŭ� 2P�T�B�aP1:�S"@۠n���5/릅rD#^Sa�����J��ċ����tGC����ń%�Zg7!���m������2M�F�"S�z��:5��7��ǽm�NiF#����m&e�F-o-��qu}�Wx���M_vrHH�1�y bҭٞB=�����b��.ڌ�cړt3_+�}N�hEhY�h�$�W*��g��:|��k���^j�8��c���0�/��'p��M��C3�!S�+��J�#�(�zkG1�Q�xB��Hm�E�khIO�c�-�R���լf���m�\����>��s=]��'����`��U;U����ή?�~i���(L7���|1 ;�^/��E�g�p�O��8o꨺�X(Y����*�� P�?�z���E�V�҂��L����>u��։(����%%+#c���!����os��KaG$
;����u�M�����ɒ�@*S��c�˘�i��^��mtW���8�~Kq=*)�$r�$q���F�,�<Qm��O�D����O� ��0Κ{P7e9:2b�~��S�h/�¾a<�4�(��U�fRƙ|OA�cS7r��+Xu��R>��B1�4~h(㏊�yyRrF���0~RX��c�L�(<D����ol��6�½۱��&U����G�����:�	i�P�n`�����W��Z�0w�ɕ�R0������ԋ��vӁI�)Uf$��x����L�d��h�=��	��ѥ��K�����k|B�n���Im���+�H�9ئ1p�o~P�rG����F����B#�\0Kv@��f|(��Uǵ�H:!��{��2���ɪ�|�SA����}�2r��-��i�B�_
e��T<%t.R#�_��%Y�I��u��PZ�%�� ����=��t�?�n�j��s!��J��Ǭa�j0|@����<�=�3ك���r���ɩ��a���<P��q��-+�[;����h����
��t�����j���^"�PR�d���diZ���O^��L�z�^NXޞ�5>>Um��M�b&�U/�gB�v�׈������u�p��X����<�X�4IrW�bb���J����T75	f��x����53�B��h�c+�N{���cC���-��ص�\&_�9²Z3N�1��~��A�N�ӧO./4��9���cc9��v3߅�J�o�N7���re�|�t�u7�um����8��:z��[K�<wI���e���K��rD��fv�Y�03�:�b��SP���'���u�iG��= �G�~A���8Ƿj�CuTU��'���m�N&ܟX��Z9v�с$):3��d�s�6��$I#?�?��]�>���ߨL�Wײ�S+|�n�۵D;3<e	�8=���GDBͫ�nE*�c"w~f���lT���}]��D��4G���+�uf�6��:�������.d�����j[���;������c>���,.fAe$Ń�����6ϔ(�ʥx<�?vs������,	 6 �R�g��B�?�J��m;J�j����ōG��FUm��]dx�8��W������f
�V��P�w��u�b�qGP�7�=<�+T��H��ίG�'FB�b�ފ�ۚ�M��f(!Ǳ�?��쥤��U[�^h(V_�G�G% �?9y~II5o�>�J&W�<[�ccc���ܙIN���nz}��n������/៊���(��,%.�%�P�}�P[{�f�A��_����RRW�մ������4�x����p��~}���Ծ�Nz�[��e���=$or�Z��N&'[�Xh6�L�!��D.sd 
.�&��*�)ccE�����F��~4�e,}�x�\�20�t��B�f�<'���G�>{�5�ړ=h(N8B�ɸ��'᨞��V'�!�[�����R�Jt���/�r2�+�����&�<�)��D��|0]4 gjT�ֶ$�����Y�0_]�3��$��$�?��Т���- ��@}�F�u-�-vF��ʚ�n*݋o6��U�O��p��%Ѫ�Z92�{��'��-�^?�Ǎ0}64Ð��˜���2\�;�?p���"�-�&&&,���J�װ�]p���J���>���A�Z���S1��R��Me�館4������ 5�#ZK�߳�{��� O����t3Z���`����ju�8�����q`�;�.+�Nr9`�����r�0"]��!��y:mҒ���BA}�q(�̿h�D���~�}=��Uo������E�Lj�K0�2�{0'�1
�G6�e�a�b��n%�^W.��=HLNN޿��w���y.��\��-%ؙ���:c2T�4�~���`����u���(-gy��Hz8��r}��(^$��c�d�l|����oky�VW8/�o���~JA��^�\> Y�
֒��v�ڑC{_�5�rٿJެ�e���&�u�V9n�����v�ceu5�c�%e�����ˣ	�y��A/P��Ō�#?��hN��G�;sGm���� !�}S����������saBN��<d�Q���{�o�A`j�~��h���B@@`}s�w<R�(NR��w�����xy�9�M��#hj2W�����{�{���?��) ��~����a?-ud5x�o��3Ivǹ���K��5fe�0��)Ǥ�B��A�	l�Cm]��f��oB����S�Ǹ������g+P9uo����ļmq�=5���޲㌣?J�>�%%�P��d�3`m�&�S��5{�����V��"A�vU*jk?���J"NEB�~12hu`DTY=���F��CRN��eC�&�$Y�S���mm�����=X8��<�0�3W���X�
>_�ݳ�s[,�w
��@0������ث�e��v}(r> ӳݎ�� ����F��2�r����P�����&SC�}y3jy4�h�~f�'>ઈ��ENC~�TF�2�r�]�����ӽt
�C��p2n�Z����@�ä��$���UϷ]#�{6��Z-�p��+��KX6�	�	�p୭H-�_Y�f�:��a�J�d������?磀'���D�����T	#�������8-�J�:m��:N׶���܁����W�U�i�e��E���:M����?���*���!��V�I=���VvSSh+�Ϯ��	0�H�S���{���9���SQ]�e)z�0��5���lg�ˉ���	2��6Mu怭6�E2��4��c�BJ^�~�a��f�Roj�aKޠ��*��/���M������,��x!����9�{~�� ���p\�WݬJ�Z�x�f����É�LQ��kd�3�71�����K�l�N��P�BhGF��X�\ҋ�~'б��2��EB��_r|E�Y�W��#�0�����^Aq]~��5�d�hǧGT)��m��������s&1lx���<�d6ڐi��h�t[��C6 ����	k�|4,c����+	7'��x47j-�y
n���8�"t�%��0���
,���Z�L�X��vz��u(���\���q���g{ˀQ�*=����������^2��5������sv�k�ܶ�]��ܯ����зڷ�;���&����!���ʑ����Gl����ʰ�k�\B�%��y��+�jj�P�R�rM�l{8ƣ��5��~����]��|���v~�n9�k`T�����`�}���*�O%q�(�.�z���ߟ�O�1�e�u?�
�ݩ���� \��b����`3�l^圈؈�%�W�t�_?�d�>�w��������h��s�-�ɼ����	�P���s�ig
�=��ˤ�(��S�'���l�Ar��7r^�l7����ѽEù�	Y�;ѿ��BP��HND?�n�y�ɮa���X,����Ƴ�	b�VvY��ᢹ`\U���o��'�k*'_�ɗ���H4�9y�wY��r���K�u��Db�zX������ݻ�h����&������[��:Y�e�D`_�b��M�K�0����_ǋ��L�
HH�w����"��:osLY��/쏞$#܈HJ��3�<�z(T�5DL��Ie[x�v�&�x2�8���s��J���yyP��z � S-}�I��EI�U�e���{[�:+�׆��V��W���&��,Yw*W�ṠJÓG?�h#�ĕ��A�r�&\�d�dڪ������ o6K��~6���K+�$�P�[��W���<1����X �K�o�w��*���*v�����8�S�(ZJ��Cq8��o��~!}��H����-�Fhn��֣1E��G̓OdP.[��Ժ������������}N����ꂪ*��q�Յ 	%��rF%�`]t��蔡�ў��J �?+EQH�%w�L�q�'�)�9�%M�Q��d]B�8�:�9l�uY�:���o9iV�a�3�T7!>��&G���g�j���(�9`k�?@��%)o_���=�NV��s�o�|K }�,�`C����lc���x@�C�h<׿�˅M"�l�z�2ɹ������)K�u�76~�҈�kT`A[��&��[[}�ǡ��>^O��'(�eߣC�eX1��w�7ӣ?%IRyw�?��%��sQ7�Q$�ht�Ӵ<>����#�����]��p�n>�����"��vގ�n�ԍ?<-�����̫���":D��F�4�����J@T�$�)����"i���%�L���$O/���ᛤ	ֲ���._��n����Q�%ȷ�����]�~��b����_��ղ�e-I��t��,��~�9�W,u.�{�9'�\O��>̷I��?��ke��}u���_j<H�qT�6
��>�C����^'萴K�a��0O�Ϋmń<�9�H
�4�zU�ʶ�J�����H�y41������)/���6���o�N]/��h�8�B��9^}m�a_2x�F��N�
)w�pdQQQ���������
�\Ff2~>n&v�I��a�C�=[u�7�3��Qo/�	��]��?|�-�cX>n�U�1�c wL�TXc^c����X5V [?��	����\�,VɌO4ҫ��h:���3��C��
&�F_6�����O��0(�g���H�ݮo����ڴNz�<֯WbCJsr�}���/�����@���+{��n�.�:(�	�M�~#QQ�9����ϧ�$��V����x�g�E�^[��M�<)r�?(�wZ0{�s`�G�PcyW��	`����.n+2��C���$i�w�r�D��7���3���#6v�<,%�z%bz�ֹz>�ny	�%OM�1ߵ���J��X�᷑��y�d���i7J�J"�8r�(A�e%z�� �t�t��c��dq!&�BͅQ3��������Q���YIcU��|�H����e�Rc�ӗ�'n;*�/�G��Γa��k��-�:VV�/]����)�$���������j�c(�j{�z�g[?�_XX�������I�ˍ����,\^6�I��{]�U����h�d�3�%A���U+����c.���k�%�����^#�̗L��]
X:%P/�u�G�?\�ݵn{]K���s�c��{̲φ�E���.�����;X(�Z:D�=��3��I�L�r��]ԥ��Pߛh��ҔV.y��q�:���ڭt[
i?�
�W~v�; n��)ϫj�%�ĉ���I���$/�5�'������n����m�F{��POBuu�Yk|� Ql������W��Q���i����t�c�H�F�J��;��$K�!�"�EJ��妛[ x�ё#X�Xg�b����Ԕ��qx_��V�"������K�SҰ���F$=j�qY�NfQ����� ��8-��;��[0�-�l��,�R��̲L�@��>j�R���c?*mQ���#p�߯AϞ0��H\Y�k���_4=0�@t
�z�M�px��^y:Qux'�La���{�8Tj#�\D9B�耹�98�l��q([	�~������c
��FEk�~�Bc�^9���>��i�,� u�}�����A��ô�Z�q�{
9@�fB�+�b�-{��n��`2�?�K��S^����H�9�	��`�]@$�p��p�T��t[�$�Q2[�٩�`�B��
m�#�t}�<��/��o�5�X����a�s)?�i�
����g���2{�i��zT?���08����d��y-�ԋG���@.���u��,sG�a�G�������V���:~�1������X����e`��<��	���@3��R�յr �y/��y�XHb"QeE��� �0�rG�$�ϭv���Y�|`������TfNw�r'����,��G��Ρ���MW2Rr�����G�u��l_����j1���e�Z��T]����t>z^T�0Tqh^T[�3))	#Y�H:w�W�A���Lɯ_���E�������#^�X������ⲥ��Cs��7�`����$�/q���غ+���Y�qε�J�,ĺ��q0;N��y���`�� �}��S/�`�K��U)��+�i�׭��l�9��5EO�d����W�<�{�zu��n'���A�Ļ��]�I>���>�ʵ��"w���B��b�o	ah)�YAhKM�H�PV��u"����"2rl�vC��X�w	��/���qh(��ȓO!!8���sAt�za9V�I�!�i��6����Nua=۩gy�~������'�ڞ1�,��X���1$���!��uo6Ԛ�b֭E��y��҆Vل�at(���朣Sj�;ZFE�{M��.%�H�<i��{�S��<R�ؔM��]q��\�E�\ta�_B�/�\�-O:�F�-\^��kYzU�[lI� �7|-�iZ����RdT�4j����	ͯzyU��J^)� L#+SSZ�����\I�Ѡ�^���ia�/9'+k��?*��xsr�9_��H.��x6/� C�g	9߇�Hc�8i�� F&3�}\˳��2���t��ȋX���l�d�I��e��ȝ�-����PH>;�nf8`�M��M�eΜ|���?��`8^۴�Q�Ӕ�CH� ���p��I�����v�����E���eSy��us'�	lfp�ɣ����y2G��J���_�����6�FF�
v��Sሂb� ���am�4�V�Ы��C#��^,��D2�]�A�<,��&��x:Τ_^�a�k��]�4����\�2���ܴ�Y��?��o8:��04�������*?|^�Ѻ��:e�,�,���r ���T_@D!��,@�G%����]6AB�3`c�ZO-�#08��,:�#������c�T�.����Z<���s��kC����֥PCi U��-�^�;�B��b�����e�ٸ�'�Q����]��6[��Q��,ź����6d�W�3F�T]���]���ְ��̏��6*N�fT��5H�
~�Y�[��W�L�\��
"&�b&`�v���^^�o4���(��߿�u��907�����W�(������
�ngg��6�c߿pL+�NN��-;�6K�J.b�eK�>'��G߮���o�u��[��^���6�=+�������<�^|)���j?�N��9D��a��-��������zi�1xy�d�Gɱ��Q��lV��ٖ����ؚ�~y�z�P�9����Pd���Cd�k��W��l��T�K�8�x�m�&�9�p���A;��*^��,��ҲX�$���>Ȅz8�0�ٖ2-e��RA�A��]+c�5ȥ����$y�L�iK���(X3��L�(>�`�h����~���)y��EEE�Ke�*i���+"22��v2�ttV�2�q<Uw�k�U��X9�{W��C���5�$���Jt��s�c��梯;4�c�.�����仜w��J��~[o�2�Rf�~|i���u�{�4�-���U��q�w�{֟��h��(4B�T��0TA��^)�k0�};��]��3���y��C,��m�삂�t%J\��m|���Rmm�֏�]�fݪ4��پ�(T���5���YR���ln7/_�s��y:
��*&X�\��j&�HF!��+�؜�r��`(���ϩ:\��ٝS��C%�y.+.�U�m����.��Q��A�/C�c���D���ySc7�s{�KW���!����ŏ!�ێ��N]{O��t p��zF�B�H>��3�׾a���m���;a'f�yď��X���1G�r�ix(Ǒb�$�����Fm'�S�U�\���&��WWÇ�z]'�~��Bk��|�)���p8���c�A��;��y����������ߟ���:7ȱ=x��wc��;J�0��q6/��QX�f�.���U�L�y^�7+$e;2��G�[@Eټq�4H� ���tw(H7H�K�tHwK�"�t�"�"���]�����Ι{8gٝ�����uϘɶ�E���\{�}�7�4Y���o�o�;�9��]���Gy� �B��ɭ�i�� p:	�G��Ղ��L	]�csu����MM�"�����\��^�Wb0���Ƨ)�Z�P��|g��x��o�F�9�,V�ڑ�����{��ԯ|��S<��orF{����A�+��^���SMM��S:B��)��px�M�*X���Z�TdR�����I8�kR�rL$�'j:��U+K��e�d|�}{��2,i��÷o�*�5�x򦿫6y���:\��uQ%��=��OÆ�5��]O]�����T++�U������]������UW��zZ��B ��ϗ����"c����Zb��ML�0��⣣�_��LxR�O���в�7e)�����r;$�Ǌ&�����i�2=+>֞:9;������#Z���  \�d��'�n�����u+�����N����G)����������z�����P�u{�<e�9�Q���NMܼn�R��m+M��M��a���"n�z��x��Fa��F,ӂ�����D��M���#�Oƪ�E>�F9����4�j��Q&�u�Tk&�ͫئ����T�N���Vk=Ѱ_RR�jP³L<L�ə�"={�E �K�{�"0a�=���n�5`�LMԎ}����2=�~��@F���x ��\ӵ׵�w��ATE��� �%�Fֈ{�B)�?W*;���K�V���/�6��M����SN.ZԿ(t֦�L��]�E8s�[�iH����]b{�kH2:
�m$��I�foZUJ�h�Ij���G3����K��M5�Q��yٲ� �Ju��e4[���",#J�x���vc1{@�6�ʜܲ� �;���-��{f�-R¥�[/�L�]d����|���[�:����02�Ҥ߼W�r~��[����U f�
1z����F_�֫!�=J�-=!G��u����Ϻ&�	ϯ���TÉ��'��!OW[���}p�A� ��	䲠�M����c\B��ť�����a��z�7�3�[qC�/�D��R(�x�:�$s����tx�Ջ}�(d�B��d���q���8���ʭe�������u�v]]lS�m&7<���W@I5ߟ��W�'��Σz(z<eR-�|����)��\�<��������������ޮ(o���[�)u���cqy{�����=t���l��9$0����5��WR��3G~S���Ho�{�LpK�b��Ȩ:z�~9cE����*���ɿU��Ըc�Z����7SJs�_�GӢ6��n,�O��!�N#�ɘ�.�!�e��?[4$���9;]����M!x��~��X�Os��`�5F>�Kz��'�e�^Ђ�Tc����x���Oy���mf�S�2��ܟԒ�����3�4@�Gɱ[�$f���ϒ��ۂ
��"��[-\	���\�~Ϯx�R][����o_�� +r���1��_���*;��la����{Gr#[�Q"�����vѥ��h6�����#|w���"'ǲW��,������ �Xd�V&&�kڟ>�e*�V��������K��J��XM�yg�ۨ|������B�Q����Յ����~WW�f�x��/R�gL�lYF�X���'�'E�p=�*�W>c���fs�{�&#?��$Q��N�Z~嫝���N����k�֐︕z����T�8LhV˲a��]�_
k%�vB�Uz��
:���,p+7J|sx��t�� �ַ�1/�sǽP���sU��������[��O�j��_I���]a��=Le}�gN�?L�T+RCdrg�y�������_��Ԓ�H����VT(�
�E�ک���lq� 	1���ַ���w]t�V�!E���p���8d�~���������Q�:�<�l�����enn���"U���z�!:&f��[Hy9��V�X���d��(((t@��c�~�����p7��a%��Z�MS8ꦭ���z��H���:4�imS���W�o@��0�}�qwuq�N��O��	*���i�
X��+a�	�1C�.f�3�,����?��ba��L�]��T�z^�Z�����"*� p�{j*��@��T�5><�Z�0��q�( �
��^�}�����w��4��-n[������xDRo�\���|��*S��L� �9<��e�X��s֢Y#G2�]"�R����f�k�z��ב6�Z�Q^P��I����װg<c(E<��f� ���]�����f�8�k{�B5��>�j_��vfQ�@u �,L�a�'Kv/R���p���q�HYۮ���ͥ0����7�ګ���LݎV|�{�;T*99�x
���i>�!s��H%�~(��iJ�/<k�V�e����MX��.r9���G����֮D�_��͵��+m���A��&��k7�M�벏�B�� �ʣȷ��DO�{�U��	n�׎�ɝ�l�ií5��,~|Vũp���ם$�����������[WL���_k���L͵[��O[l5�2�Gs܊�����S*@\v��ŴQ�D��Q9��,]ڈ�F�����xȥ���K�l�Ҩ�����G8�1:?~`o�w2<�?�{��W���N�ͶKۑ��N�Q�1��7�3't��^S0�Y�
��[��-��ބ����"��f����i�QJa>�h��P���I����v1gљťҵ�G��1�����?<E���$x��}N�-dn��'Уۻ煌�m�~��?����΀��u�~�������l�h���K,��`X}.&!E}Gd|�Z22���O�>w��#�Sg�Oj��l�Tppu\/��^���\�q|�z�^�$j��sI�O8��ށ�Nv�tb�<�O+�u�6�+�.���>���?�lM�\vJT0���Kl��mg<%yS�TaV���w���@���ˁ�ҵpip�; �?owkhY�bf��kh���N�Rl`)Y�i*����eo~^���GŌ� ��E^,�UU-�Ga�ށH��%��t�b#���U�����{#Y+I>�֤]ta%�T���9�tr#���3e�D���Z~C`3X^ET����a��F�:���� ���zd7<����6���ԛa*m��k�|�Uz�Ӽӂ�|!�A������YvwZ$�uw��L�C��yC�ի���k2���=��i��m�͙t��3��;K7#�N:[,MC\�؇\�d�j��/Hd�>.T��^���f��Ȩb``���������0`�c���@`=�>^V��y>�-�\0�-�)ɲ�I0��9��$-$��ejxz�_�����w;�c1aG:l�zT�?�����-?����S�S�xΩ�Kn�(����y}�¼�:��{�gHhf���:&�
|J�釣,�FN���CL�ﶆƇ��*R��nw�۪���r��]�BԊ1�2���A��?�*uO_��L�_�2���a��lU�ҟݒ;���k��u~�ʪ��a��ɗO�Ƌ��(Q("��_��n�H�P���lL0���,rA@�8�2�P�7ӰcN�RM&
k���.w��Jc5b �Յi0�K��v�e��0y��"z�ud�8͇��>�]e8��T���=�;obf�$�R7x����c;EMd�C�q�T�v�Hz�,��X���p�ZׂR�����)C�n����բ�֬3�j���Y�w��^���T�l���'w�t�����ǵ쯇j(e~{��im��+���@h��/3T�IIH��z�"N��U�9'�KS7Q�Z8�<�^�
�յٳG�|Zy�f�4��z���!�s�`�w=b;E�-���?�8J���������kz�д��[��A������piH}�t�3~������	��5>O�^u:O��]�Fx���U��$b�,3YJ�,�_��[:�ߣ��ݮ���R�k�A
�ܭ�eCp^8	}N�������MMX�Iz?a<	mK����+�-�t�r�%I$P��2q��ڡ^af��$1��L9$�K�N�5 �9U�VeU�m��O<�����o��a�
P9ac��{�~`"U�R署��0!h~qR"��#�~����V�.S�\�r����b����O��%1�@�oUUx���"W��U �,��=GG	j��yk�qMމQ��9E��k$3--�?��{	�E�h���i��$G���� =Y�)sp�}�H�����x�]���K9���q$�߽�����GO��M��JkR~b�}���i���t� �V��̘%���?��6$>�D��6�������j�� r؟y�� 2�#�*"P�9���G��v+��B��؇Ł OU��(����N���c�Z��*����P,�="_>>�f�;�8^K�?���]&2���0���NQZDo�z�N}4z|���;��$�j]�S��~Z�MO~o�j��q=�Š%e�.v�X���0��~������,#�.i�/�*]rK�Y�Zy�G��}=��cf�7�o���А��4*<�c�1^�d� ��wq�k�����+ה�qg�Z^�YQZc
p�'�d�
�hQ����ػ mˆ@fj,qΙ�7/<i��-E9G�:�c�?�)��÷�a:ޘN�١�\��g���=h��f�قV
�>ڃx�h;|n�S+XlA�M�qT�M�����ݑ��W���i��18p�Ә���͘j�[z���e�?�|�cy��j��Q�uj����WF����ă�@�,0���&���S1-�Ϻ��{���a�O�����!�h9ҿ�Z)��ـ'*�����4dv���k���h	��x�e�Ǚv�n��n=2&������A��f-���~[�\���d����?�[�߄�#fe�R�������-h;Ƚ�o��/A���"��~p'L �fL��&�H���@����gv�*����CP��/ם��>/8tam�7gZs��	猦ډg2}�R�@����/����p��(1lj���}�Դ�F�Wh�M�P?�Xy296j�!;6�h�A����U�n�Ջc�FG����|�wf����5Ͷ�ca��n�>.҄^������7�6���Է��Än���j��]�FM�6�X�:Ժ�s�A�Q#zBBC��
�`Q��D�jX��[8�kM*++� ������P ���W�lZNEOxB���(�Q	��;�t7�sR�2k.�Ӯ폂܊\�35�A�[]i\���5�~ch�J�h��̠��D;GqѨ��A�N�Nw�c�zSPh��d]�t��O�Oǹ+VX�m�>�����a�铻/
��؄�?��B�H�3^5s���q+,zW�a.cڤ�]�>�Ƙ�n�鹈�H��tQ�O�7Ci\�|�.�IIIK�zqey鳙V���ҸHh&��V��@"���愤�������N<��5���ɒ�'�o��f�@CB &&���I� _�;�Ķ�嬤�X�2vG�/���E���3y��.[ޗ��/�ڒ���,:�S����`>\�,e�~��aa�l�X�~%��Ĳ�H���ܮ�=��vz�N�VVV������K�g�ܼ��>D N-δ/]�)�zcK�z|5�$�G-jdL�����H�e_���E��#|h:<��O�:��Z&����j[��[��8^����E����,�Ê��[Ea8lW����k1�X��h�󛶥�M^�[���#��:�g�Z/����7���޴�Tk>-��������T�>�r���}�%�_�\�Ч��r�LI�_=>>ZS��������c���28�g�Ib�Ј�Z����\�����,�����v6o��L��bF�d�Fv����j̜�k"O���z��q���Y��@"#o<����C��yy��{{M���KQ��^���{	3��m^�f6�$�u�*O�ﾚ�(���o�g�T��M@�s� �E�������8g`�݊_tz��R7���J��OJ�+���a�9�������U�&��ƭo�h"�Hj\�94���"�هP�X�#��^TTG���:;]Q\�������$��J-i�W���݋P*��{p =`�T���gu�������~t��:�7��Gz<�NB���cY�.����w�rvWlEֶ��Tf�lw���J����~+-!e�sVl\�FĔ��M��z�Lm%]����^�YLU�%�e�e)@!!�.�lV���9�]`��+���y�y�j��_��=j�뽠���e���xx�E��|�y��x�������j�K�����$�,���"���O�v(k2���ۈӈt����<|�r�� ƺ��B�2��G~,��|�v4���$�0oߎ%��)�!{��_%@G�w��(p)�5�H>�����O�~��U�����:ɿ����؃�8�bw��R��]�=Q@�N�?��S�J{_�%,�{�yOƫ$ؐkK"\R.y��R�x�6O��>�.t�H%�5d�ϡQ=�ss��%�><iu�}����YJ�����`��r�y��O�tJ$�v�r��8�,���6�WȠ��w[�6�7��6������#:�`q]`�ND3��e SWͶM/�W�h"x�U��$ �n0]�����������+g7��/J���j�"��>0��pĽx��ɋ�`���0K\\ ��Hj�����'4����|�g��ʚ~rlaJrQob�		)eOA[��xvd͐^������6�6�O^k_$Z���-jv�ʹ%�4lĴ`�5�{���?��tMeEK�PD>=f����c�<��2` ��8c�r��'�.'���#g)�����Y����F)ܱ�&t^��]��0څ�)	��b34}����.����gb����`�P�/��D�����7n����P�@I����Ns���e�؇u��W��\cI�~3d/�����Z-D���@�¼X��T�#��#YB��?�Kh��.p����nE�f�M�"R~�-��P�Yt�)*�[G��:�R~�	-���[#A~u����̜�6�:�����T~�$);w��p춠��X�˪�I�TK�9������g�qW)�{�K^�%QϮzc�)����w�Oʘ�$	���	�q��桡ܸ��^DˎON+f�v��޿K0��*V?	��ڞ�.:�2����:Rs�:,�,����B�3P�]iiSS��n�ᦽ1�J%��u�z:��N��퍕��R�?L�=�_D�+��a��~�zS����KR1{:���[ڴJ�y�9���BD�pp��%^ԑ���Ͷ�����!7��l�x�t7A������?��ц_��L���(���%��-����������lU;:����7�BJM����hU��޵cOh# \ �|Ê��w��'��Q��Nҁ�KYB�i��a�^���fl_�����^BCC*VG���� ?��E��T����B9�M��]��~J�������{�n�bu��f#����Z��o��|�t��$x��왽=�m9>U'�Ѿ^�j��4-�U�����^����nl��<�U��rd���.�}V�Wy���&9k���K�+K����Q��&�'�����gK�?n�q����@$x�a�g��?h�������qI7+B�J*�Gk��>�E��<Z���F���.B7�$�9p[�X�v�	?��^�Q�򥣴n��G\��Y��;T�6Cć	�kS�Vچt�A���L�K���G� �kC=y�Ҕ�&�#^��KI!��9o<髠�Ɍ}4�]��7n62�Y��~��2S���n�y./|� �1`ط"&܍b~�7�i��D���c���%�����e�غ8?/�9����<S�t�R�j!e��'�#�
ITS�L݉��Z^�I�S�'�7��Ȼ��"I��5�
�ف��E'j���u��c�	c�t�����&�ol�� �@N#c��LB\3T��|����D�����A�(�7l�x1�յ�2�f��Nh���ZP�^�5�U-�ʞ����y�k�*;B���NGS�
�Ю1W��h}6�i�i�ơ��6t@X�>�Up`e;Uک��	�F�N�[1l�O��O�l�{b��;�tB荈�gr���}?��Ղ�K��):k��4��E����O��b�",�s�)<Ї��^!d���=�Y�P�c�v�)E�.�q�Q�>�]�������jJ?0�3�+I�Z˽�I-Y���ngx�@���g�"��dW�Q��5(n���A�o�d��(C��_/�Og�dg"#�Ƅ4��<�i<�ͥ��j�Z��	�Hq[�ϊƻ�]!D&���d'9�����e{�مմS<�e���<i���ߠs������D߼��_8�>w�49�����gU�-�L+���F����<I�Tǧ��@�y������Y�A��,�~�^����M�vf~n����z��-�w|C�˽M
yG�ߍW�`���8��C��gf~kߝ�ZeA@����
+PV!��O�q�_��ު>�u��X���g:�����y]ϚB��D���-.t;g"�-���!bf��m:N�B�j�mצ���L���Y���5]�n�'�8ł
�g��f�gp>>>ڵV���ŏ?�kL��y ��G<���cD��Di�s��*�Ol�ZԯO�,)Ը6Q�U{W*	���)��`��*;�s0��W.<���aV-((p��ۻ��7_#[/q9�Y3�YH�SaJc����Y�怨X:��)i�
�Ɔ��>�pL��ts=��sJ��gCv���j"��({ݻ�~h��{�}iHqsy�>������nV��~��+��{T�a_̆�x�JӮf�_���,�}!�)�R�h�7H��V�6�7#�<PX�kC.d���[JV"i�*�~�☥-d�R�oޠ�X���(�u�,[� Mb�JH�ݽarcH^Q�G�7y�S��;�Ʉ���g>�$��r�)�+�|"�1�3e����(?��Y�{�??�I��[��F�r4�; u`���A�0p�F�&�fJ�l�6 �g���u��~�mO{�Qa�S��D�~���]t�cZ��c���I<�w�@�nP�����+NrZc>�nP����r�=�x��I�=��j=�u�xSY�;���>�X<*� &B�p�y��.�Vр��7I��&����8��(Q}� ���v����t ��:��h��N� ���(��I�bfA#��j�'7�P���N��D�[ ���� C�y�q�Ix�Ȑ�xJnR>! �śڳ�ꌿL/�I{o�p{�в���e���0�v���Ne���1$��*��)�^w�N_�Rs7�E��>��o85:���~?T�ڿ�S"���ykDFK+u�\噖���J�O	������5��u|D��W����@W�|����~S+�V�_M��?�i���R]�;z�\�^��N�^�q�K"��r�tΧ����	��lX�їH�]�{���L��@�7��w���nݳL+��l|>�*d><,*�}ቶ`ta�����[C��I<�w	���5Xc<���<�_�%F-sm�-P����% �8��p�;yR��`�j>��Ɯ6O��8�j<�f	q�A���ay!��E�9�e����PM-1w+?I��������s�Ol�Զ�/�m���{<��P��O��	q�H����;Us^^���+M[�R�?�_ӜN��V�;��m8����f��ַ�1�ϓ���~}*|r>�O:dZY�~Hܘ>>2͟��5G^��v��#9��Ϛ������'��$�Ԙ�,JG-�m�a�~�^�����2�݃e�as4gPL�5)�bҷu�*ޢ�m�����>CF�s�ξ�
N:�qQ�n5����-��`K�b�	�r(����	�Ҕ��t���"���7�&�7~#��a֎i��*SX%���� 5]d�F�9Z��v���D�?�9����Dx%�����gw��f�R��2`�\�О�B��Iǎ���H{wtE�7l��^@�n}�S���������LK^�ʝ��)����P����䙻��8m�F!%Y�����0����eՍ�U���\�?^���F�YQR�kK���q�A�H���d@g�z��z�H�h�h:1FI3G�+X����
t�h{6�b�F�����sw{t�+Xhd�v�Ш�}�p�+��UڥV�}��z�ۂ�o1���ʥ�B�{�U�4�G��95釸](1$��w�Ì<g�]��nI����b��f���f���p�mX���F$Ϳ`Sy�����t[�p�40dM���J�E"��Wz	E������\�o�Nə�g,>Sd:y)�(���VO�b~��{��Phx㘀�T=�v%\�fُ������͝�5)<�Ir��+薴����!]CP(􅺔�+ŉ�`*{oO4	(���]�P6́F������u.8�����F9��/zȀ��g����p5�l�&����pɪ�%��4d�>lUP���,�w��<�|��Gr��b@:���\�ݑ��Q*��}��@��ޙ�m��9�;
�<����\�k��W�<���iZ+�ʦF���cLI5=ފM��N��=�<�Uo
n�K~\�H|MQ���P'��x)�؞�QyC����,�ט����w�������c���<iJk8�X�K.�[q��O����*𽈎��JU��m�,9���˻�>�byY�0�N��	-�3�����|��cV,T4�{���n���Л�خU��Վx:�8��J�n���ZmM�g��V����|�~^�2��ꯊ�����W.�A"�aq��q"43�eq����}b��zk�Ǭ�߯�����A����Wwm�#�1u�N��>�㋓�y�k�_��|�[~�-�9p��'���mA������Kt�lE����)h����S��V�Z=�^7�Ӡ!S�������TŒl_x�24f�L��\}�� .�#'�%4�dI�/8���d��@|/Xu��gl]ڽ"���Ɖ���;��p���s��R-�J����&�缾�wS�
W��e6J�������=�w����hk�?S�*�k�]�Z2�pK������-�ul8����Ƌs���{��T�t]������o��Z�긚�'�����,�i
Ps�e�.b�doN�m��SZ5�d�O�0��%�!�>��eR�dlv����mB������M�qL�ܿ�,�7</���Лp�}�N���8�\,z~t���e��yߚ�4G6^�"�[�'�ָF n���hk
9͎R�~'�����Ŷ�u��%�������)M �����d��-�\jqS����T���+R6�&Yn��1����L�l�}l�
�l������ߘ��������>�.�o��Ã�}uxx
p�v{����`;���%qKZb�����e�@�;�R鶾�>n8 P�ʻ8�����D��m�//I�X �* q���o']�٥x�|���B�
 �H�ɗ���X�6����e}��]�3˰'��Ӗ��ΩBE8�F�_�(�M�ce�U9��#�����7�'S��ˏ(.|l|(c.ge�e�Pl:/�4�2���xb�K&]1ݥh���{%�����Em}Ո��}3�RlZp�J|*����Cii==�͡����zG�˔�����L��a^�;i�^�8zy�OO�.-�_]�>�[��~��̽��H�@���(��U��mԠ8.���~�g��-�;g�=�W���9�]�-��:j�h�I����m� #���c?��nK�\�N��<�'l4���ID������ܒ�b[��!�1}n�ٕ\��	8��n	�>���\��lo�,��A���E������� ڧ֖�^5��9�������OQ���}á�%����c3r�x�U�In���s[Qz�w0Y}q�碴Y�����/|4��������R،�h4�=@�a�n����U,�h�ۏ�����~[j����2x�F�Tvn�M�v��D{��"����DK�AC|8YYY���?�S���?�˞)¬�f�@`���^ 1����S�mlG$����)�>�(�F�W/�>
�[V%��@����h�s!��ᇯ��'�a$G,6�Q\Xh��aśhN���"adD$Q���N��3U޾UJZ��Z�,��R`{�V�^^N�@��������;;׬��abaFcac�.y'�h5�L���c���:bu�c�Mx�����~�IC;K�r[t9�J���(`��+�S��@��i���skc��Fv���}g�~�JD�u�%���'��F����.5-Ĳ�KLCy�u3[*�'	v�x"k'd��%Q�jӠ4�j��O�q��
f_�[f��D8d�?b�3u��\1�Qn���$�r��Fy�}w�i�(���8���y��D�'�\� �\���\J|�L		�g�T��:Y[��	u�A�����斖*�Uɡ1*����&�b��Oo��]:�,�����擲���L'H���EP�"�ot�5#=�����Ԩ�׎0�0$��dQ��ȓ��<W������x\ny�8l�&�hdv+����Dc�r�e�
��L:���5:����yyd���	�b�������q�<�A	A��o�G:�W�2�d4E^�7p�ʴ�nT������٥c;/����"��]54��ꁎ�/��/h\�%�s�����?�W?0�i�U���	�0��8Գ�34~Ƚ�� $f�?����c_��V\��Ǎ��N������ �f[�L����m�6)e�����]&گ ���-u�dK�.����_,������Y�칏�-������T�f~@�K�-���c��%x�f�!�e�<+C-�6Sc�u��)U��t9�t��4����[g7����\�Uh�]ͬ]����k�^�}o�gsqw�ki!�k !;�:���ׁmԄ�P����[��7�ayUUx��O�����&�zc�|����I��ǘ[}m'ݩ��6jt���^:V�4�T� ��0�3��ݧ�u�`��\�h����.MSkA�T" 
�)26��(R��ǈpC("-*�3h����ՙ��l�iqѴ�5.2����s>˷��X�#3��@#N�%I�dJD�+���� �U �>���Y5F�A�SaZ%�h�;D���0��Z�Q�K9u?�k(���ʨ�f��P}v��Q�	k�|�6�������#Z��ؗ�^_���0�����c�F��D�u���xzT�ً����$y�"���7����vU��MNjLaOB ������W�����h�ՙ5�E3�Q
'��v��"-�K�w�ĆS��(`D�'����W`Wm �:�H�,�;�``��Zo.���,K���\�di�d���r � ~�C�nB��nF�sss�l�$�P
8T�Ȟ�,�X���Ԅ��8�K6��Ⱦ6S4����Xu n~�O��rl~rl��?�"'':i�Q��l3�\9g~��+�:XX��0(=\�`�K�q���M�� ^�1}�Z\��
fӄ�P��S�B�.��=���U�8I֒n�r�ґYBo��N��=@e&���i�{.8�Dm��抰E<bF�(���=���䁋n;�Y��-��ba�τ�b�"�h`���w��Ld��֎�F�����-z��l�R�B��I��d�
�Pd���s�ZA!����p={(!���r����ZG �L�=�/�3�7��!!(,��h�J���{�B���ʯ�¤�	�Z/�΅��&O�+g	v��(�w|j*��vJ�@~���J�&�'���FO�n��R���i=�Ȃc���<�iŶ�r��E��� �(\S�R�].���|$�\�����Z�x`>�����E�n	��~�!�d4��|Ohu󇍡&�}�?K�Yf�`ۃR�����	�z�˼ܛu�I&�K�?^~��s�Y{��hmuZ]u�d��VV���C�H�Bn�`*4���¸�D��A� )d-�=��6Q���)<�YK���$��n�YuS����))�1Wg븑��c�L�_kve#�D�Wf�i�g5�p*�˓&j��R��X;.���	߫*[7${k�ٻ4�����2=&��m މ�o'+�&&�v��v�N�u.�qs���ꇣ]�V����0���e��=��b�5���VVLG�4�DsB!���2hUR���ӈ������542_l��������1��l��7�@���R�+�����ʸHܼ��/"����lmaxP�VbӨφ$��h2 c�Ud.��!�?�~�!���78��+KK����1'}�������Ss�S�p7��k`���`)�k�J�;h�(�j�G�x�e����e�X�P�����ѯb��@8��~�0��nBX�$�f���L����O:�m��8�r�$���c*/���o�\#��m�NJ��ֲ�
�������W�·��=Ӝ��1n,DRc2��� �������5d8Ӥ�I��O�вx�	~�!�f`��*�����(��B�P����J�QJr��`#)������|U�Ю����g_Q�*���0��H^{<F ��^��5��f�D,)Np��Ԡ�a����n��W���ë�G�N�P��qݒ�S#�[a-M�J�,��Q��<�v-�O��L1��yv�TXe;��
@-���$��n�*�@���0���`OP��(�/�%��}���F{e��7Y����kҗ�4h���d�8Q�7�����R�����Gc4�υ&ma�\���o�����q���\&X���
�'iӈC��:,,������"�{z�����L�+ƿg�݇�o��L!�~Ǝw����>�4���%ڏ�	-�Iǀ+oQ�˔��#���������&�ca�4y��t���;�?�W~�����?[��u�߹����*����)����̓[�wFp�ӿ��j��=�qT�I�E���k�Y^t%�T�-
�(2���+ݚ��+�f�C���Xx���,����vx�W��Ayzo��O� �%���چ���\����#&R���"�m܁�K;W����]}�9_j>�O���i����
�to�!�:T����IZp�_ǎ߆++6,8�}�;����=�����g�n�#i�}�4�"i!d��|=R���(0��'��TI-q�xؼ�0���Q�z�d.�+�|��c�H��T��!�"êj���#;���W��A^:���e��-��zΙ�	4��i�HII�-��N���8��mf�ˊ��f�xU�?�0z\!2�'�[	x/������{>}r勲6����t�r�{�EFEB�Ks�󬐨�~z� �z�Y�W�ŀ��m?1>nkkK0�J��[��;��Ǯv �Z[�&o�,1-G�5kd��ǋ�{�skn-�p�:O��f׽��m>O�2�~����N���l�=N�4^Aޫo���&	@T�qBP5��`�Oa��0�/Mv�9W���}��>�шh���>��F�!	!���������s�aBP�at̪��ls�e�O���2=�[z�7�T���q�N��Q{�� P�}n��bH$��n9M�ǔ�[L �ۻ;���������7G�/�z/��b�*�)���a݃�W�
��߼�	�O�>m��ue[�C���3���Y�����]\�m��x_0���r�ָ�5�I�,�)bK��0~]"�e�~��5��׿�Ѵf޳�ߋb� �AB����)¢a�W�|(		�]!���t��3�+7�U�!�� Y�.°����S���BjZ��(�7 ��v`Z���V�?I�w��'I��ֈ�=�/�v��K��Gb0�[4�F���t�p%N�kM=t�p̫��Z	\���A��E � >�
z�3����˴R�����&oA*�ccp�X�lw����CU�i
�\i��v��) �=�O��F��19�ϕj�\N��nM�Q��t��|���z��Z آ/�)N~`���J�{l�ɡ����畦�3s��?�|���.�A����-��4��X�Ҧ���v����3�J�a���EM���8���8I+�g��Y��^��N�C]�	���ThJp7�"�\:H��	�ѷ�WU�����w���!��(&&�d�Z��ٹ��˅(�H�܍	�Tcb�I���O
�l�aE�Q�*ue�t��_�X������:z�Zo��m����/�yB�o�I\J����!ʰJ��֒AjYD�����~	܏�`
���Uߐ�Bi�R�&|�6
�"�~׭ؠZ�[�ȧyu[�7��ء[˪� ��L7,S�)�!Lq�,hh�f<�*��.��� ��m6�p��#�D���n��Q9����H0��G��I]LZEZN��fD��8�͖���S�v#�in,�׼��c�@|��a�oĵ�.�kNjf��ΰ�v�А�����l�|^_���u�������ea/�|d_z�̮�*�chW�>���133���o����xc3l�
ņ������͘�e�Y�@��o�yf(��.W�����ʆ�m���j���/��.'p~��[�+��B��L��%�\3z�-�r~�(S���&M7E��[��|�B��?�3����,�����7G���^dN�/}c�3f��Z03���}��u�����v�q3x?��԰�Y�YY0���ͤj&J� ;�2֒�l�p
��Vvv�^vV�!f��)��.���@�<՞y�20 b7��$Z�ʹ��]r[r�[|�#���<�-F���҆�o^4n�Ko��u\��������6�&Y��D��j�J��l�ֶ|ww�֣�Az�*�?����M)<v��g�'��d�}����[D&�F>^^p]!@�o�Л��I�ߺ�� ���%�NK�;׬��E	! ܲWm���
�*����/ݍ" �)� ��"��Ҡ(H]����D��A���;/���1w�q_߻g���ٳg��5�T�g{݈�ϟ��:�Z(��jU�T���)��߂��WJA�0먉83'��'�Odv��u�~���-_V����Q��ܙ3U?�xy�[�
��k7�������!�5���f����Xy����I'E<�WW۽𶴆���G�A��1WWY9��gm�h�:t�����.�"hRFٿs�����ď�f����s�v��)gc�B~�5�eH/��p� �'œ���� z3^��
�h1';��;n=|K!�J���Z��ݧ�5����1�o�S�f��{Wҁ��	a�Q��6��p��m��HM�S]9%%��SV�c��Ʃ�#�h�����z��)�̬���X��q*.�<O�<��������
�a,�0�3�t_�[?�X_j֛��5�g�����K�k��qO44K��$��NE�П��-u�_�D!��[��$�'w��=F��;Ư�F���A�՘ ��	g�IZX�}{֕�ض�� Ha^��X1müX�z}����7s�X3�'O��0��t�^V2���T���MR�O4@�zA����i-�U2������_�9��v�z_s4���Z�^W�	a� ��,.�zJ�Ȼ�)xT��,�J#g(!� � 5��db�>@����, D9I�����O:[��.�n.j.�����*-�uRw��X��p$~��i��$�n����������t��i����	�����.�
Y{�Z~�`k������R�=#����� �ڭ��|�?�1�`����;}�d��St��̳Z$;��t��唜-�����]e:��Ч��ӓ�����[�P1��&�PE�f\Q�e~�l�H����3>�a]e�F$�|�Gq!�y���Ne��bD�j�8�l�$�hW#7:�Gm��Pބ���̵'L/t=�)��;g���>t�})�c�]��E�6"qCΫs�U��ϯ���ï�ő�Y-	�Ǐ>�),��p3����.���ֺ�/}+�!Ұp���B]��x=`	�f�e�	���B�i0��ˀU��9�6_0�v�fg����ؽ�2�VR�-�?�s���i���T��v�}�����Ϳ�B��``���D)�yA��<,_������M�Kꥎ�5�J���=��W�Ax����&�XyKA�qn�o����#��D��j��A�t�j�Yy��c����|��$i�ae�G�� �� ��� t�V~0é�1��tL�'z��H-�F��Uu���΍���~�aאˌ)�Z�+�=��w�ҡuv�qa�]�~ w�7����4�]��V��U�}�I(k�F�����}�uT� �D���=�����ā��^F�3�����8���[��E���Ʊ��tHt�O�~7
^M�!��� ����h�u!�h��P_��:nM�����v��E�W���H`xG�쩻hף�1z�����YYL��+$:X1�t�#+�!]4�g��}[h@��V�g	�h�-֏4�X��z��y��L�PU,!!��֙DPx��
 ���E�Ǻ����!�NNvwS,���?��P�X��-�ڕ~����є�� �[��qzͤ݁�����A@9M)i3�o+��.%%�K8����Bw���ȁdӂm-tJ�)��P]�ǀ��F���Y�	��_�)!G��\�a�-����9k$�zQP�I����@X�`,I�3�w�F<tz����bɨ�QS��Q�\j�ܼ��hR��n~#�p�	Ob�>Q��^��	;�S�0K�S䖎9r��X"!%�뿋��������Puk����`Dp�1�����m��F�4���,?��޻
S�w|�M�`�p�-De��b����%`�^^b`Q|[��O�3��{޹s�t��3�*��B8/����a������&�&rҪ�|M�.�{������,�GB�/���-��<�Ѫn9���5l� �gff���S-�8tj^�\�|��v�!��i�G��ܐ7a�����p�ef��L)�՗�$E�gϰ�u��mz�� '����SL1I0�M�G՟Ϭ#�����b����G^�$��uQn���fswFj�f`����lƉq\��1�Je�̸�]m�i����8�0�F(t����H�љM��1�5u��IW���#�{�fo�O����p���#��Wl���x�1T7�l{``�Ǵ��Bk��o�tf0�i.��`~  ��>h����6��*r��U}��QXXx:�"�]{�z�q�_��՞k�sa���2�����/����@�� !3�L��p{��f-+���D�Z<�]#��jr�y�驩�2/i�;LL�D;�57�/�m#�h�Sa�KHL�]֑�2w�/�� ����Z\��I�W�7ݰ�hӟ��~�*H���8�OɿA�hP_��k|����g,�N�)U�MI�ە��*ܛ96��/��B��d������%TU���W��uՅ��ST
aď�)aI4p
Y���v�߂��9Q�i�#�+6=�V�:`K�;a!�?׳ޗO��no[Ae����i�	�6����ĝ��&��������M_P�V\���n��yyy��}K����D�}�~�����P��{��^@#h�l&�������;廉�E�pݫ��`׮J-,�]�5'h1�(VI{�2�ూU��#f�3a���S}�Q�tl(mc�f���`MS"�>�~5�e=�@Ks���=����j���KQR�A�uW��4ך�R�n�{�=9$O�|soϋh}Ua�ޏlBe������99������#��4>Y���z�L�������%��)�eE����9�iшl$̒�'mW��|��̡tW���\�2�t��ns{Z^����٥��k���Oũ�{��\�Ə��L�h��r�?3Ĺc�Ԅ%/���`�F��= �4��r�x��t�H#�U�H7B;��̺=ڮY�(�=PM���L��>����Ђ^I���|�ߒ�a�3�A����ڵ@G�W���К��z�E��׵���;:K|��~i���d��E���b��ۭ���*S^}�Z0�������guRRXS'k.cc���8�z}� k�%����v(�ڍ2�d���&��m�e��P�R�vq[3�N��ԋ3�3!��8u5�É�6�4��n� z�}G�a֒��yc1_.nJ�V��C�o"�S���7f;�ӧ�\�5�4L	������A&g�~Ρ��*����Z�ٜ�Zu��+\4��b�Nc�F������ޙ�|�����R�1�3sԤ��1K�1E��+֊�����C�w.΄c,}G�9jJ��(qN�ւ`TUS[�u�i����T������[�#����0:�!(ck[�7��<cy�з�̯��N��qOO�徔��i�գ��K��$,�=	�����ә� �Gߣ�q2h��R�6�HÝ|�/�/�,�a w=���H�A���;m�|�#$K.æQB�����0��"��#�;�Շ�_~��I�h�R�|��̋>�"&Ts���'��̣@�F��\�[��a�[��冕Z����.�8͵��R	���:�6�J����frC8���P�~��Q��ɘӴ׹;L��>�b�s����feϗ袕$�����w�׼��x���Hf���ˉϷMJ%y�"'\�X2�^�B��
���{�Z	6t�A�>c�\�3W{���+r2�GnU�,##��6���f�;/QQYٲ�r^^8�6 �SSF���Z20�e�������}�L����'Q�ݙ���r�:�k���<�������-��~���JK3�ѭ����E^���GL�^���+k�$��i;��a� �Ԋ
8S��1�K~����n�%�+����[��s�-�]���d}�F?����hi����\YW7<4�I5�KLl��o�A3 �%��q_Y�P2K6��h�'Fk�l�{�dl��� &����秈�?l���mL��;�]?��2���4�J�Hܩ��A�cu�p���������I�Eo�+T�s�-���%���\}�cag�1�}$dt;*����V���)|4���˚��2�b��-޸�8$�c�b��<y�o��+��Q���B��F�k�w�m�<��T�O�>u���P��5�#''�����@�ʊ���@��p�Ǧ]�F�9Da0OGIG7�G�]�G�f���bDf���g@������5ϲ��[�4v�&?<	�Y<k��g(�u���MXF3et���W<����%�����>)|����Lã��]g�����T̰��8]�t�T��\�	%e�b�G��V��P�E�M�@ Jn�.a���w.�{�4'yS�AB������W�K�?�ؕ�R]ܾ�x��r���8HF�g����IX���g��W�N
��e^��)Q�lQr�����k��c��CS�6?ڴ���U�+B���E.je.R�M'9���^@�F1��l��`z
!��8�oLL��z8�V�qӆ��^��� ����CJJ�2���UV^�707	���+�������*���G�{����%44ځ1>ٞq�-�?>N���wQ�U��>~oX���Q���c�I��?������喝��I�QjԞ�B�0j�Ǐ`�8����K�t�ӊ�����~f�� �e������qK ����|��|r���?D��O��Th�[��b"ʔԬ���˽���y��L�d�wOr02���eB����3S�L]����Hj��˻:�����Ҍa��%���6�S�5p��X��D��ê�5�K��F욋��B�&��'g�S���J����'T�����{�Ԭ�b�)��o��
B��b{S5�2ql�gi),�Q-,���P��[Mr{������b���+yy>�ԑ��ߑ�W3cE!h������)A���eM�{�C��B�p	�A����^A��w96Y�Ⱦ87�k?�]w#4-*1]]�>�E|�JC���So~���{�^����Z= t��L��<�'���Y��ﴏϿի���(�\J����,�L�U�9������?T�K
)�C^�`M��Ϧ ;J(á����5?�r��yXo�7!d�!**T���%�'�LHv�Z�d�sՇ��Ž���3�C+OB���	4oL�����g����3��uW��̹���?Ny�z>�LO'��M~�.:xN�U�H�M�1�N��'�Z|�s�ovl��o�"�χ��$�%x-i-5#�f�'r�'�$�b��������o�����oGJRDB^��àr!`�SũV�'k��ЙŪ��3����x�4�Z�-X7���({��)�`+�`�Z���N��K��E�K��ǚ��(�*!5�e�D��xQy]m��c���䊖~<j�CG'x/|��E�����˴ՙު��!����G����5��O{����Ѵ
�>��~����%����s�.�����̃_i��jz���l�)Nc>����s_�F�NH �:4����+��P3230<�!`�!�Od(V�*W��oGݶ���(HeKJ����6ڟ�zV��&OJ���0���m��z�-.����g4���ǎ����i+�[ ���H��Қ�|(�Ց��.4V�:>.n>����5 ��H����y��l��	KYGG�0�ƻ�l��>���X|usSآf�QZ��_@@���3���p�Y�Ռ��~=��r����t�Ջpi��W)�a�N��ncsLa�"�p!���uH5�K>��z,��������C���,����M�s�����%�c:U�nB/~x��~_"Ǥ��N��h��+���ȠF���r�~�jH0$+���@q��YW,��{��*�lS�P[�K�g̊��PH�7�[�!������~7Կ��ύOB�,����*�������	4��v�JD��d���~`fF�[�Ck��r��y�$�ֵ:�����S[ɇv?��ao߽�NN���'�hUw�'�'�?;;���G�����F>�}7��hhh i��-[����	5�=�3 �F�6���>�#,,�9	���v�L��A���J�(����1g���F��:a5j��?�����(/��B�&����r!&J�
��y�wNJ<.�k������e�o�������h.U�uJ���wK�8,-8�?������	 W���MM���y��Ӭ�R�ڴ�۷o�'&\��̡ҵ�������CWLL̗zz����k.���Ձ���\	u��Ӄ#�>��M�G�{g}^�I�!������G����Ñ��S�y�z~q� ��ۑ��S��,�%���=_���1���fN]��kw!ܯCƨ޼�|v�F�-��o	���5�v/�_ݵ���V���)�ac�����5{N���a��m����v:�L{J5�Dw2|\ѧ�%�*��Ü��CThT�^ ���`��D1���U�1X�O���^U�|����f�[p�`�qd�P��xx)���T��>zU���K���h|��knβ��b ���\�ؐRT�-x�&Ku���/�ܥ��-���N��7H��I7[�h3����n�j4y6$��� ����`���m��r�ׯ��� ��S+	ߓ'�Ӱ�]'�8�<���@
�@>Q�_�A����G.����jU>Q⸥�ܠ�9^z�G��#�ѽz�
>�S�x �4�;?�������b�w{�n�U1}xN�V����	��a�K�;@�N���72��DB�8��G���d��%[��e�
�T���@�]]Ǧ�y��8 : Βn�����Ӹ`@x��GD�:'��GD@��:�����FFƚ��B{�MW8J�g��>���o0����1�]�_�᥊��c����lM`�N�
���Q����M^�w �O��"'(*++��QQ���M�Z�Գ�$?�=�z?a�I�ug;���I"?��3��r"����#Wh��G	`��y�����t=\���dddP��)^]9�y����_�9ƪyg���?K�m=����?�%�=��E��(_opV�3x��G�ϭW:�C�u<��|=��| ���z*���J>�ɛAH,�{LZ����eT�>[�����w��9�����B�°�y�t�[�4�������6E߂�YV�>r�sJߋfm�h��� �ST����B	���]NE�+�/�-%��^Wb���;0G������̌�R_�i����Xm.���j��ni?)	w;�c�����<G��pa�|N^����yI%%��+�	�,�%S[�VN�Ɛ���=�2r32��yB��Rϝ$T���f����aI�����eH$��j�:>z�]N��Bֶ%-OCغðУ�]��g]D��1}BBN5����}\|<�w�GiلeHJVV<	]��w� ~�VU����;��zs���|���,�<��Qutա��R�K�D���%�j/z��=��W/6�AE�oM�w�	b9 ��O'	)�4b����$��F�j�/�R3R�O��ÖԞ�f��v=w����\�M�uc�8��H��LHϴt4�/Rbo�쬞�DZ��N�O9��_(��$�t����N�5y�Gc+���e�'���҉�ЂBN��$)�p�\���`�x��m]Z,hck�=M*���m�a���3*%O~��1A���t����P,|�Y8��PF[�dYi��-�»�w �K|�g!�+3�A�%g8(D�FqS�8M��Z4������||�Ư怣�R�RTn�� o�5����MM}���X�y_�֟��^�-�H�锁�x?o'ۭU��������߿�Vd ק��ze��� Rκn�����>�U��[aҤ y�/�Qe���Ҩu焎�P��ǹ��L4�ė�'jpF�މ��x�M��q��h��tu�/v��s0w�� N��EP|=��S��SY���C��Q�-��||�E*���j��a��0��Hˍ6K�PIE�RRZ�G
P �972_&��ѡ!��9O�<��3w�$�/6ˡ���O�i"���������d��Lq#�\9��b(s ��+�� 3#���X:��7yrtl:@d*�72��P%>Y�s�c��!�n|�̸����4_#5��4�U�+��=Y��.M�g$�]Ao�4�&��_��0!�ƦC䚢�>.x���>P���9��D����Ϥa�;����ϳ����O=A*Ey�E�6��Q@JrtHߗ����4C®��Xg�W����}�m�w�5̫� /+�7d�0����KE~��_�wL���	 9JO/g?�����sW~
\�7o���[�����cs2��(�$�p~��K�?^.�ZקK%� �� X�2��
��S�z#
�ѓ3�����	��v��GO�M��Ձ���S�˛C�եS
}�97&���J�{5nR���W��W=��hW�bs�Omv.)WR��v��w���A�V����B\\6ߐOV���*���e���>��&h�;�����S�s6�i�вN��L!]S��@hj���'#W�Ѐ�r��q�?6�B�'���RF�ݠ&�e�ѭ���Ӕ���=���U��v�ٍ��qq ����ޡ��&��/���F{=,;�[[%�]V�N/W��R����]��7�g��TS�v��;s�c�TΚ���n��P8`yM^7�8'�������W'sr�h��J�?H�4a��eU��Ed0�(k�ZW0PQ��jDի�*�
s��:��-�9��2��5��}l�f�@�huk+i�I��u|��J��I��xER���T�JI�̎�F	1ƕZ���r�ʴ�ܡĮUi����G ���#i{V���>Fď�_��1�{���m�8]]�Uh���s�֛!&�����:��89���YB�~����x�ص@\��N�		h�NkQʘ����� |����8���OU�`��M���W�k�k��.� ,�U����ee1Y~ol�*��7���6��FKZ�P����բ0֏t��O�g�pT�����(�ƀ��.�	�ĪP+�)E��U<[��9��m��<�k���kg�1�q�vS^I�r-���3��DSP[QsSٞԨ����XF�#��)�y��G���Ma���ש�4����BG����%egg_��	�t����fE���*�C�� k��SS����or.�{�5�|���8���?q095e��Dk���x]�m����*P]]]�[Z~;>KOO���?��	��y�/J�C-��[�1g�󡶝8U�`��e'I�4E��(I��}]�.kЪ����Oq�c���������g���܄�,'|��%���2�3<�}#��a��R_���I�e�n��8]0܊���ö����4�F����!��tK\�0p�c�$���;�6{�VqRRR ��3p+��!��aV����7���x%�ܾ//T�֠��l9����������DI�ﾗ��P�h�D��U~0��	�CiN���>�Ϟ��7R�#�G�q�#(�
-@��6���%�_o�Xw��w#@#�ۭ#�� �&�ߜ��ӧ�8O9e(N\ӫ_l�l�{�I�JL�	
����>B)�{�ȟ%UB�Sttt�L�&x�%�G�w���X����^���Ĥ%���Hg?��V]B�^(�SB�"�u[�P�4(	_&��q��m���y�'�4�|�٨u=K(T���qk1�W�WTW����l�t����*�Y>Q �.�C�UH$##���${�ZXI���n���v xП�g���L�d�����D�r�MοVF����KW����fT:?m�0c%�wCy] �RYYY&*l�R���;�f���#1���̟�]�ޗƱ�h��-�|�{j��x'z�����2|�ݏ��Xh���-d��_�Bxe�(�p��L
8���������;��ܗ��C���fD����k�
4?C�K��Im��`������ ������>-Ï��f��#X��#��#Lp��_[�� �9ӢJ4��� %lQ-�MY����lmm�Y7�%�m[ �CH�P�'����p�\O��7�8��A����=J��vz=v�ڀ��Qn�\M)��';r�$�BY,��Y̴��c/�eM{u=��r*S���/w%�x��?����'�x7hK�n�>�2c:���������a�γ��%�ł{�V���(����GAW;�}��̛��)��?#��g$Q�Q�|n�n1`�~�z�P|ͽ�vR��,�%y���4dd�:�y�}f�D��x�_����ujE������ �ml��s(F3܃�]�H�'�U��Eb������@���ݷ�2<�������2�t���i`��7b��jj6�d �]hb��8?o��uT9�2�7k1���"�$ l��E���4��A�\ �^&���g��_3"���?NA��q�6q.��]R$l�Ψԁf���1�0{v��^��<�صC:���$��E����u$7,�DB*�ŕ�S-
V�)���q���\�*JJJs+����Ϧ5:��%a1�YO��m,S�*c	��8�G
�&'S��_T�����!$�H�L��q���%��	�N�GB����p)���O��̀S�^U�HH����v-j�VvW�w��V�-��N��q�����*���<��O�4�i����ލ���e6">Y���3>����,�_}�6��i=;�7��o���e��t͢'M�qy8�2�Kmq�ts�Q|+���,��o��]��9���������`E	��)S�������A���f8X��&i��w�Xo+Y88 a������2)t�	���iz�z"
h���J�8݋&NB���� �>��Ihkk�XY���s�zG�o�o؞e��n�G���p�$䴸�N0�w�9�<��A��������l�T'��)L	�I�*k�����T�h1�l~���|�E7��ۭ��vE�kb��x���Nݦ-`���(�\Z����ص�Z�"*<͇�J%Q��لݗe߇B��a���Y�>44)B$6��0|\G.�0�R;ne�}i杚.(]���"z��Nf��5]r!�Bۢ�.�:��z u(����5�K��w^y��mU��N6�no{6Q�.�455���	_>��[���N��
U��4ݡ��ݠ���[r?�W�w�HGO�P6��~����X�n2Y��.뗗���T���a�.A�w0�CT��o��ıoQ�����e=�0x�����L��G�P�
Oۖ1�m��� 
:�A��EB� )D��0��ChBƱ���}?鿿o�#����6V��{�i�@0���_cY&� YH�"�������B=r(���;)����/�L�gb�zY7�� ���@�=�(N��D��d	Yل-�能=O��f��DW��_
0�Nǭɀ�m��s�W�,��,/M��ܙ_�B�����JV���1%�d�K����NNN�Bs�)�j�MTFR��ߣy����UWΣ"H�+���=�Mj�W�Qiؕ���|}���)-��ʂWՠ.���^�F��i�]�H�;	�3nkg�� 5b��EH�A�\��V�K?��H۵�H��v�~��q��?R��O��ښO�A��׹�����CUi�8�
�Λ��4����t�tCɛ������r)i���L��H�{�� o�|\q��?���~R��鋤��1������ mP/�H�T"��- G?5.g����q/෬��o � �7�!���%`�?�|�ص ;09�h����0�r�4-ㇶ\�M��IRz���Wl��I�?o�p�k�Cϗ�ME5��K�6��%��}�'??ߦ���ْ��"\�2 ��ޝ��&���t>]�ߦ)b������	���8w�]!*�@��Z�E)Z�equjG��0c>Z��%�C#��O£����B;Һ�3�{P�V�Jr[JU5́o�_�=�����Z��Tl�Eڃ'���*q�"+��pqe�{�F6z��{�Ώ6lk�����=�Q�����k����Vb�MǕ�A��̣e��E��M��2��W�,h�A�Wz���"o��������r����r19�R���
#�#��F�$���)4��vb��wE��1-G��*"*%g;�$Š����¯�Y����MW[:�ܨ�>�Z��9;m׮,f%Z�tq ��0y�:�ˋ}�����y��O��ƉaRT{֋��I��To�o�V/٧9�nF|����;����B�8�����x882	�����v([|Ѡ� c=QĽ��'�CK:���i�9?%�y廯�$�D�7%l��W��l�JH���|��J��8�	��@��x�C�;�<�>l��H�,-�^�k&j�����s0ʷ>���/���9���eb��U�(4�쥈o��a}+m}b����K�0�t��쭈ݐ�"�3�+,�sq���@v)����ާԠ;c�:��d��4H3}�D�Py�K~���ǒ �%j@�FR9�oN���7�F���COA�&�˗���n�~Q���ݘggg�mi��0+�zL4�,I������T�6��ۻ�U�[4�"k�/lY<�^��Yu_����hQX�SS �xr���%���%�D�F�mPJ�-Y}y�e�o�p����)�P<c�	Vub�ٴm{NQ�uA�)�;�-!8�@�8:��p�$��%6�R��A�~�����4a�"�p%�=�KO1�[�_^�ʃ�j�����9̞ˑ�䃽Nj㡬 �B��o����Es��v���,�$�������<|ͨ���r�Ho7>���3�Ϧ_z�st���ix�����Bs~q�	�S����5q+���3I�?��.��N�8�F#��Y>�v�.���ܗ�Ӣ�/��R�����1�E��Z �'�
�{T%���_���g� �U��w^��` � A�-Qd���1��/^VV6�L�TE�>��!��Nyp����c~~����;�>}z�*/-�sbf�S��$#�f/c����h�#��y׀�5�d	dt���7�����"���!X����.W�m�M�,�:�S�tg�z{:eȒa�{�=�^�v���2��Jwm��0�����X}�BA4��b"�F!�-�İx�
͇Vڳ��h$7X�Z�H��$����	
_�n)А��iEii�������fO>�����A�2B���kH�22 ж���8!��2�^(/�����5؈��<���r��z�\!&�]����<�*N�@5L5���[ �}�,�o�p�ma�p�糿�mDy/2���!�4����h'��k�����M��Ԧ�����!cQ�L���O|�$F;�1��"��Ux�Ɩv�B�c�@!�ЁZ����q���CY����s�Y�Cj9���Él:(�O��ѾM��e��&�������#���#��b���_���E�^��i_A)���.R�o��eNi�Pt�G<�aۖ��&+�XX���������^3) �L4_�)�)���#yj����!PDh؜�y!����>����Iv�R�Y���������g7w}Ij���[�=j�K�$%%e�E0�,�f=��:���񢍇"���w�Q��X}iXj�oj��NXL7� ;��X�p��f��k��7=���]�v(>��Y�Z���%������G��߭���Sp"	���ug5,�W��?m5�h�;C]d���<���ք4����|j~�^�5
<�qV
@�p�\#jIn�#/�o�H�cf0ڛC2��� Z�ߓ�	����U0���_�G�y��O��|��;�'nН�� ���6#bB�2�>�3���X>fw�]1tGV�)阮�h�f��Lh7W�vN���J������7�bUU����PQ������3����]�¯�=����ɩ�iN�����ᖌ_=w��ώz�"x�s�|H�VK���,>lły[�:>>��y4�����@�Aw��2��*�4��Iw��<̂��]=�,�9��{	�Y�w��{F.ݟ�4����`2qz�8���03������ʶ$X�b	z��:9R�_z@0�:!���������J��ŉ�j(	뺩�R̝s�C	|e)�h�~��pR(��İO�|���Y[[�΅��{�	��4�`t�����*�(�AU#*�K�n��������@����%��uP�|6�.��pVm)�ՠ��t�(x���h�\O3IĐ�e(9��C�L�ٳ����zL4��7��2I�l]E�嘛������y�|�.��\��A`�;�'g?n�����&�_����I�S$�̘������H�?j>��ʧ��HJJ2\=�g�a
Y搈��ʍ�MmS^7�J�����\���1o�"a�#y}�_�	2�_6�/#����E�[�?�.� V�����[I��`	eaa�p����ϛ����m�[�y�!��x|Z� 5���9[�X��:�,�?���3٠)��u�N�Z��\�T����2b A�����#���O���",�ۯ}�"�囤ǈY�jϏa�-�����͑<BQ�+m��O�	����9�#��2��Z���Ge��RC��Ň��O�	a��P�hG����vM''>��5GU�@��4�=qorZ�}������F�Gng��9N(��x������^���ǭIJ`��g�T1���[x ��t�R]8�"^<���n����w��Z����32���
���,|}�U�99BoǠ�.Cu_�kA#�IU�����qG,u����Wz�j�>&���*n�>?��s?�'3NK�^�K�R�tlӻ@��GH.=Е�I�&e�*-K��vz�=$�W�LO�M��WWb�y���b�-�)̈�B�=//Z?������I�m�$��` xi�P�oKvdm��t���	��qFH8�Uhݑ^и�Q��>����-��L%2�ĳp��´��N��]׆��⠹���b9�N���/��W;^�"n��I�Q�"BD��5�@'u^�* E�c^��ί&�É����h�z4l��m"��B����x��\JA�5�78XV�Vs���!�(�� $]j�NN:}Z%N������#�@�)'�����K+��|ݙ�����$x����������H�͜�}��oi����i�>�>R�����1���z?�(�>}Z��"�]]��뭭[D��L����@N���`��;�(������y�Ɔ�\+��.��2/v�T��BѤ�zT�O���fW�ݬ9fㄵ��v���0�D��3����qd�<P�o�݂U���L(�ʔ��*c�Ujg�z���v>$3�}30>��<4��O|Τ��9G�{DUU�`k�� �U|����p]]]åc��qi�n?ړ�8�[��qk�g$7��(��o��j1���>E\�ɿ	w����F2j�4�����m��3�
|�ۀ��"$��UҜ�|�HN�G;1��]�Md�����r냗��quS�������A�����?�z�/�W��5f@�ˁt'�x���t��"�0^�Ǳ&LGGG��ot�9������gr0�5�5;${�!�t9�˰)�&9�0�\%a42?»�w[;.no�D���ɹ�@GX�����ι�vk@��B��F5'08�ő�V����u�۲� ���B���PVx�[JY�?�s��'Wb�1�S�y'�e:96��ը��Ą��fƬ<��Y+��(&1t���]���CE���v���C�U(����ȝ跸o\��7�\����-/]�m��F����,�e���r�hp�Q�Д���;�e���}QN^?��5�@8�L�@gNȱ�}���l��eu+�2ʰ���{��.������n8 ��88-+��I���Όv�l�+9Е�ʖ��$��<� �d��0�$ۖ��c�S������h�[�y�H�vY9�S@�����N����k)�u011�fB��7�}�n���-b�zq@�z�d�k�~�^X�߆��{���3���H������%Y��]��F��[�K���fq�������%�KP2���E\����e1�f|+�E��Z���j���P��-�ׅ�������hDD(�I�1��@��a�3Zl�K����hd��-}F��'>���"f��(2j#�L�&�50�������œ�_�GHGY.�C~��}_���h�8,�+���N����^�#��P�YZ#��,�д�R�3�v�X{�N�q�?��:����^RS
�;r%����o��wN������h�M����7��_;ȗq�^��j�V����mya�`a���!C����Vj&@�fJ��\\\�O�˦�Cc� ��-��{vo�+��~w*�K9 ��v�۟��(�W���%��.�O%�dY����50@��C��E&�qq&!�A��=��gԮ�y[�8��AFQ�]�����	U�����60m�k(|4�b�G�����A�A<��r�X�/�j^�1��IH'^�C�O�z?c�,c�^"��cMF��,�j��)lQ��z?@�b|s}�a�͎T�� �m�)g8Lb�,���n��:vr�(�}�{����ô�,��G�"\\\�	O��
������L[��'� yi�K�A��@�?���6g�%b�x
��vw�m��\�㋧��bL���ݾ����8���0�	�ݽ�t�賷�3K���-88�#PeKFCC���A�Y��k���r5`sW2r��!%%�Z�����3u�Z�D|��w01[�^���}���v�NU��s�g��x�#T�;=��x��Atuue��58:�I�]=�H.
�-�W�E5u1�Kn�S�d����I���}���9���k���[�P�ޤ��>��t���ߕ���⿚���gb/v]�a��b��yh1`P�Y�^ ��T��ⶈ�-����ϊ�K��oZ�=�aZ��L��^V�e�Dz�/..ʷm	 ��j��m+�J�.Z���]_��+ t���Zz�|��ML^�y�|os�3�����,w��승��e���o���z�#����E�b|Ǆ�������Q�XG�`�7f��Wh�ubY���	X�3�4��;�O���g��pH5و�-�r�b�`����Ս��vR����>H����N�A8}_�aT�L>�'��SS�]Q��a����)�!4�VY!����y���!���ܴaY���]��Nn]]�ZF�fЗ,������7�]>Q`�	�<D�+;}~�İ�P(���N%y�5 �n'�@����d��})�x�]7
kNf�J?�5�^׾�~�Gמ�����9�x�S��T��o�]�l���d|w�^�$��*|&fy��tϞvQ~��1�PQm�ߣ^E�t��tHK��tw��t34("�)0�t� -94�1H����^���b����y�{�s�y}2�Z�ms�^0w4AHL�QUE���՚Wwl���P^^~�H-�r	�:D�R�@��|%N��� *�C���mS�����A�� ,�w��c2m�g�����N7o������ò���,�X����- �km8�y]�k�������gO�hi�#`[\���"b�7h럳y퍾��黗����-���+]]�]��m��M���{�j�����C�}+[��SY�Ι��Ϝ���?Zc,�y{X���޾x�S�Ë
�h�9U�n]��A�>�DVYYh�,��:w��=%���߿�G�0�@rlb��Ϳ�����5 gNc���������B�s�{{���(Y�����C1���!�9�A ��ɉK����^�5�Jo��#SS͓�o�i����P�1sy/+/���!bz�k�؊�/ݽ�}���+�Fl��:Ek@*���� J�}�*��$�mU��K{'��cQ�֢���P���.���&�i_�� �_g�4S
�X����8�����p�{6�^D�N�1<,,������T9�o�z��r����(����<���$���RUK�ᡡw��$��`C�J3�)��cJ�	H	ş6������f���'�H+���ΐ^^��rnT9�����".>����uyhwy#��5�'�[������E����_[X|���{�Uo�����b<��%�ՙ��O����:�i?>^�M3eѭ�!b}�P¾����nn�Y��L{���"�GR��4.�M���⟒�ƽ�IL7�n�EQ6,��UD���Zj��t���-����6==�ck���{P�۾��9Q;nF�	�l�k�P�qXO�N����TM�>0�:��Qu��!�����E�L�-����V�2���/�k>,�3�$�H�Y�����~���5/��ޞzn�{^<*����K���č�T_��s���b��5vx&hY�>B�t�+.�|q�V��M�vf����;�/�У�*�f¶&+iXYoC�\�����W�`�>�>�j�ƠH����L�i[]Rj�`�h��/Dd�G���'{�!���jñk�^�ץ�ͪ����;MF�.���i�RDf[*��(1�9�y��5)YY�������w�c�0G���`�۪�JRű�4�di_�t�	�c�&�֍���ަϦ_�2���X-c�ڵ��B�[�����}H��?0?"d#{���<��t���5�l��e:Il+�X��bt?��ܨ���^��Ds�L������)^W�c�_'���w���ձ�����m���J�û�%[:����+��'��̳���c�j�O}}E+lQ
t+��8��{��ʐJ��q�څ"�3��Уe/0gs{=���Vo�AbzM���'�A�7�����a^އ��R5ؠ�c��+���}��Y܅@�Ԕ^YEŋ�gK��!	�A ����nQ�n�xi|��8FT��F�_7	��L8��c��J��/x�}�d6�]&q�ٿU�|�u��U�@��b�M��BBcbbn���`����ҧgV8�(|�{��_�������>�.��Շ�����GBz{��j*O��F/�]�	�����������wo���ߡ�ލ��`O�DebbY
����*ъ������{s@��u�w�+�����;�僟��?Re���	^�q�q�|����e]���|��[���~,��IE��0���E�]S,���=22%MM���S�8�L[s[Ҋ�_(����.�����J���I����l��O�b�AmI()%TU�ǣX�@{ʐB�~�����z,229�7�u(��~�0(�le~&2侥p��!���5�k*/�$+�o*"?"���]!�	���WRQy�������@����?�L������z P��*r�Yŝ���T`0��m���bq�����̎�:���~q1�@+3�5������'�i���@�*')D�Bw����
J���n�m�����-�Px�py|�X�\d�;]!�$x���'C?�����b�p��5f2�D�b"�#�tX��]����e|�b�����pZ�f�(���T������0���3L�g�]�����a����ar�����Y�x�3Ӣ��ܰ�_O���qG��mZZ���p2�cE��U�U���Ó�r���	C_x�P�=RH��&6�R~��i�Y�:��ۯ�A$��~�9P,)H����L��k���]I��^��'5�	=�������X D6�x��s�Ҟ%��D:�ë)B��$$$�/T��-F��#�L�4R�!����Ѽ�������|5�)��}����1S�K��h>�/��H�����:d|��f�b>83�x�����̬��F:4��� ��P��Ʀ�� ���۫пTWk�џ��"��!2��t{�Q��J�b����?�9=�j��p�-��6KO�b��):�[��>z����N�	�Q���)?^1ʔ���XGd�KRWQy(�)���g�a`�ê�EnW��(r��*}F2)�`f1U0�4 �Px�i��[6�3m/��K��� t?�>Ya��E|��qq`�MMLXY�)���
��o���J�_�;iJR��ϋ��@h뛛jpxeMm���t!��iQ]]]uC�"��Ng��?8�rf�7�����unO�zɮ�WM�2��=��^"�N!�bd�|����k5��d�<�
I�6�IG��R�?��{�}]_��;Z���c5.V�
X�(D�����?��σ��l):�2�&T=ڪ� B��:!͈��щ�i�f���ɂ�\&W��^����{�]K��t0#��/2N��}�V�L||��r_��əut��
>S��n�1R@Df��%�0hV�1�?π���P�vS`����I�����3�Dyee��W�u3�܏|��f��[��Z�܀ݻۡЩ�D��z��icfb�Ty��q��9?~)�ٽq`���P��uī�_�|7�lϫ���q륳Z�9)���ۈP��3���o%m���h�iqj3R��Άݵ ���� |�����$+@��g8�Q���U�\����c��Qwy���Ht�{}�6H����=�Тmt��n{ز�P(�.�����	����\Κ/x�W����}��|���S�U/w�,��n5�Â�<2g�RI�w� ��ڢ��Q�����,����S���8��Xuʠ^�u�R16� �P�3o=Q��=rM;y�����%�s�s^h���h۞bim��\i��.;XP9�+B����%$$�^�����R�F�����bx������Q�� ��>����Us7��g�=���Ū�k
�D�����1.�'�Jj�SO�����y%�tU2j�;t9�t1FT��y��,���50��
Li�_����*�N�\dOT�V�U����Qt,7�7_d�󩇷����̶:;ܒ^�_��355�̼��������Q�����z�B"�����`xw�j�����8����쬈>E���.A�5����-:::��_��M�lUL���L��dq���	� �4u����N���>��� ��,��2 �QN}§E���!�Wa0�w$ab���V��=��L3����պ(��!}O�t2��|�B�z/�K�C�L����e�a�R��>-��3vm��Ѿ2{e���nO.��SR�r��!O�A�����bG�KQ>��2�x^�x<j���p&�,�n|�%v��5��~������1�7`�[0V0�d��?���������p�ә�m_g��$���A��q}�O�!��JJ�G=�{���F��0�tv�|u����E�g�k=|3e�t0�{��ޏ��N��x��/j��'�t0��'����EF��2>�%�3"���,�����$,�FX�7���JlW�����C��kF&iPV���ѽ��ֺ��Tac�}}o倴('G�ǧ!��i���#  ���V�o)�>�.�8N	 ��v)^")��8��ibAC@��	�E�;�a��O����q.��v�Aäʒe�sJ�d	���%���\�?�����8xr�.�]������B�3��p��j��{��-(Pם����ܗ��8X�L�m���C����Fn�֎�f\]�Eտ�Ю�����D�7�:�(�v=v�d�F~uS�~�_�A���#��uk��1M��L�n�:����u��c���[���܁$=
��;/[�c�n���a9Zk�iu>?v���yd�B�f[��4r�����OH(Z�Z�0s����w-/m�K��T��fi��g��B���k-��j����� 3���h=�VB�w�d$�П��/'^�M�IMY�ܛ����A ���y��+w`�!������1��|v^�l-��X�|ζN��Rٽ�d?��[���8"ǧ���<cI�O.�8hZʾ�O�����������8�S�?q2KI��x����fPV]C#(�������8�㜳+����t�e�v��K3J
���̽�~��4���4�IP����*I,�<��~�t5з�BT6�����=���@���V����Z��ޓ�1�ꇋ|�y_��j\��#���a��È~`"+l���$--=�{�ʽޠ@��y1����g�pD����?Ж�vSqʙ�V"�����>[B3*Η[Z�ǳĞ�0_."�ˏZ��HCӲN�Ҽ�@<��B�B�eD06:��lZ&��Hx�ǽ��
.3���aԢ�	�5� U��!1fă=��AR��E�S'�d�`j�����F���{p�����~��f��s��M��mo�m }�f_�߳ �Zk*/J�b�ު����?گ��[�S�����dt�K��r<��5�`�&IRRr�jtC��˴�N�Ѿ��~����v���~�}U�E䨺�s�H�xS�a��T�ZU^�
_x)tӻ��|T%éԹ��'U����+5q�$0�}o�b8W���E����x�S6$B=CV���L^�-��خt�:��\\\������+�i�2�HB���zD5�� ���֮��8c����%A�B�b��T"׈�q��UQh�c3ei�ങ�.0��r344�^w&����u���[-C?j�I�,���h����l�4�?�SQ_m^�K2Q�:�=����{��e�qT���,�_�S��l�:_��V�����(+ۺ>L�r#��b��(7W���jp���9�Cv�(zőhM8���!x7�M��`c��(� �[cq"��	�����[9p�/�R4A�Z��>�`cc/��`��%áU���Rpd�<��@��t�ϟr!� �¾]��槑|��5R����|�Y��3"�e[i����"r�yTJJ�z�������N���B`0�us,����g!��Mj��u<����̬����ю���d��OK+��AY���qk��`z�A\�W�9{N�����ard�i-��Vt8��n�N� {�xgAZ_PXX�˼7�s5:""M��^�v�s��KT�!.��s��}Qh=m����Eej	��-�2h��*�����:�ؕ� ��։Rs��-�,Mw	`�5�����F�b��9ԫ,y��Q��^}L��ᑑ��%.NNn�Sg���!��k���3u@5����K��4�󊺎�/,�̚b��QZ���^��;��D���oř'��Z�JUSU� s��ꏃ{M����A�ĕLp��5�M \�£Pb!�]?#���:�I�B6dע�5�l+A�������N�=#,¼��A?�U66�1�k����ׯ^����4F�t�0s�U�k�Si�TgPtq�w95��R%�*7�K��`�r�|m��`�o�*�Ǻ��4�@�� ��L��2�ܧ�a���B�Z�v"�S?Dϒ�T����_q���ZT�y�È��yy��3w����'�z0:�wO
�ԥhͲ�A��4ӟp��;���*]�׳PY��ny3j �A�DR=����2���b�V�ά�<M�e{zz�Q�"�� �.�=��	e���������y���DII	��e������xl��:�.vN�ݡ֐�9�T�Z�����r�=��ֻ,�_�f[=F[?������\K!v@d���A�/6ӝ2���,�N��H�wF����q0��Œ7C�ڴ��_P��=+�#B� ��u��Om+'A>���<v;金H�����>��|NN���p������D��X�O�<���◵>�g�P�{��Keoܓ,������ �����2�����gĒ�D�r=�y���t��f�[�ow�u �c(Һ࠮�~�u���y�=���hy٬�x>�>ܸ���Xj^Q���7R��R�(�{�vD�I���nQZL�X[1D�9�6���CJQQS[�T_�#xY�j��U�*��ط�MI8���vf�e���A�w�T���55:R�&��<�S�!��l��p^U�^ I���;B��{֠��]�'
�|��-�rt��"c��(�����I%���YY�No0/�Zit�1D!��zL~_�����[SuY\��~��o�㿠�y~�r[]_]URUU�v{����jXd�-J ����3d���üx�vi���ޏ��x/�^���Cft��}(d�����~3;�������ؖkO��'O��dD����K��9.Ɍo����᮹o�텹����&rY�=�]�5�R1��/	5]�ښ(/�����ߤ�;�tut|� �����؜��}FϪJKU=7(�Si�x �@2���C/�rS�}�vUs>\����ƕ,E
y���5�6�wȜ)����&�Y@h�yX�`.�D5�jj�����K��u�z�$����N�}���s� �0�M?wbbbz4Y9T���p�ָ5Yy4~�������Z9����65��VM��M��ܗ��l��SDX��+6��Z_=�/��ս$#��4k�^� vP����Q0�@iD��n��k�QT��H��ά��fo</��9��Kr;jٕ��v�Sm��A�4\�=�$4
c܄66�78���^���;[�~�J����\+1��2:g�ZE�l�,�� b�~ v��q�W��\Ӑ��&�O���2�'���5�F��Exb��E�Dk^�D{/7�}R8��i�ˬ�+���G�r_J����|�
��_C���G�h��(���Uy���K�%=W���A���P�[��:	��rtttL���6";n�p��5=���-��x������Q�=EB΄�5�c�2�,\`h���V|�D
��`�[񌞤d��C�I�@���@B��:n'J�	�*~��7'#ø�x��p�]mCԟ���>ꋤ(§� ���<���} {be �K�,����ͥ��O��.K.. ɏ?�$����B�x��v��})�{UZf�=����F__��):ķoJPw�nȯՐ$u�_��}��^�.Lx����#jY���U� Q�w[KA!L�*< Hs�����\}��V�h�H���3 ��%G�DH�7٧7Q�4�)3 #NI�K�FU�^	  h�nk{P�� �K�U��SPg��TPh*��g������٦5F��q4��+)��X��+>�H�prR��yfhiiY��t;0J/^����6b�j3��H���[c�'�T�Sa�ڌ�n����F2,SY;�՛�������c��G�EbAx�������E��G�	�����n�k�R�ɶ���]���;����%�W�-�ٽk� �rۿ�CFc_l)�N�c�����VJ ��|���<�8��x��X rCc��0˂IXUr���x��]�;rM}m%%�<�����i���� ��F p������Gp�4�q�����qk^��FQ4�`�9��c�t����eW�)��\���4�=��������^;��-J2��:{{G$��3�8-k�,N#��>G���.��Q�;BiM�����+Ip&��}4�5I 0,
�a�ĵ�mw�j�N�ҵVb�! �S잩���7�[��-����-d1Y��Æ�wRt�
}��D����C�QZ����~7��%��z��u�GR�j=07�zB��i�	���	��6�@{�S0�+������S
�gׁ���t�+��� ��z�����݄�ֆzѠ��j!t ��J�a/���VZ�L��o`�7�8���y�v���[A&>q�6�����v���٣3�CkDg���N&"2���aecA�d8��^�S�ˌٷ�����-�@|��0T{������`W2
t+m������j� Z����${o#��}��ؗ�YH��#G���������K����(�S̷�v�Y_2k㌝EL�#��K�z�O��#_���q��s3"���=��Q%$$��K�[+#rbl�v!���?Œ�Z��� cRR�z�R_��XbN�\�쬬TMM���h��R~C�*�'�����#�T���wD/r�C;���-�$C���LC#����T'WAWn��/u7hե�%::���켭�.�#M������Z�����Ɨ�>==>�8<t������5��,���-u�hE���M�iM���_��c^� 1��UK��v���9iii3^ �+�fD�b��u���F߯�X:�O�)����		y ����"��[!��}ް�4m{�ڤ�+��եK똾���o�n}o��p�f�rFH@���AZ 8 ��0�����WN9���6l�w�^G�e����o\��5�I�9>�S��8L�j�(��%#'g��Ǒҗ��K�s[D�7�h4O:���|+��|�Mӓ�n�R0M �V����7:�S��}�i$F�ݻ�����hsH�RO�7j�)HN���NJѴrf���
�tI��VE'�K���:�[{%�*�6	�@�#��\����tx�v����ABX�+ /� �Xn�������W��MWw7y��́���K����S�:U�i>|�2��q�vY��d �	J�١�8Q{�cg��<�^�w�`
vP"\,�\[8>���90��rn�j5��?�B�A�5'�	��VOy6쳽A�t)��K��Hŵ���ƍk�ӌ��,���?�� �G���$u���|���		�	=f.��9�U���dCkKk�lfaaaF+pi�f��O�nYO�XK)3�K~�����X��`�]�
�ݿ������N���)��vϫ��L �y�K�T�f �f1RVMI�������۫����Ѫ�/�$Z���ā�j�ۓ���(6���QI�~�۲��)l5�BHDԵ�Ki�8���q:5�2!��
�9Fn}�������Oe���{�򤴷����oa�0�M���4HĻ�D�,��J�EdgK��Q"o�M�@�6ۺ���q���=$��~�PLK����n<.F�"7��~=�5V,rF5@,0�e��茢g&�F i�%�h}h�`¯���$�L$����i���O�����g��q�pV��FY�������F�G��'l>�s��	d�ff���7a���� ������6b\�/��:) ����A�.窥ބtt��-~̒�Jl.ϖ��jq���p�)aI��ǔBnJ�L���(�]Qu���76]Ӑ�����n����0�1��5�8Ӧ�Y`��D������ţ3S����'x=_�A��BTԿ���:bV%ElF]�s#�j�5z��Hi���ϯ+��0^tI��Q		V6��2j���>�r`����m5��t*�A|?���<W�㓬Ivs�b��p�����]��)vrV2�<��u>����9����,yU��3��j�oo7M�P��
 ���5����tx�� 
�ܽ���Y���8�yu����W IݡFsQ�Yڷ^��,���3�����(d^ƕ���L�s d}s�3-��9{�Dl�'&H��!A� KOn[�:�<���2z�`D�y!G�.�ͧ�M���P�'<Y�W���Yz��ḣ"O�2�Q6@���*�,���j�m5
}e�a��􁜇R�3��Zvw��d[[5v���8n��&(*�i�ϗ��>����-(����=�Ȯ=��?+ʝ)�z��/�U�.���O0>�����������@���: 2�9dѣ�s���������>�h��s�Ky�+/&>�����}~|V��{.�Є���S��u-:�S��]7!IRe�p �>R�X�3'}�%<�m\�9���H*#UV�o+�����Ԣ
+*x����p��}/={� ;��A�\ �>��F�2�H�����/�?��׊"�I"i��R_Hb�7�'�ܻ�ڝ�p�#4J����N�cWggg�	{����e���������"Fۿ�aMW]k��F򕽽���AM^���a�{�R:�Ž�	b�Dh�IIyϊ4؅Od����X�qa��
�˃1�!Jx�����D�iP�*�"�C_��*oMU���ʦ��7�����S�!��r��$�@�A��U-����Tp}0�OcS+j��ؾ��K�����-��b�o��I�"{�}�f�;��4�H�:�ѭ���*q�G�H�9�(�8;g�?�������u+��A�o�aݟ��[�W|XF���_K�t>S�$�Q]kC��j�<�l0��~ ��;�Jߣ�T�o-�;C����� ���M&|^�����3E�!_L_����Ȭ��޵��3����� �	�F%���{�Û�t�q!���3c���*������TZ:��br>0��*$���'�5Y���~���B�$�YY��P`3i�^vE�Idu[�D��#5r��k٩bX��x艉�Wآr��c���xЫ��	 q�+��WZ�Կ m�Qy>�j���y$�&�c����i�����cia���ނ�����GAZh�=���_c��ۍ�Е��7�/Z�:�D�yc���I���E5�bW���Q����	=s5"Y�D������JVV��.�� .�0F��,��Lq� ����Q�B�F�"0�����S����7Pl�b-9`$u����^7O�uM​|��6.d�!�֮ϡ�&{!3�[*}y����N���5w.`��2i����d� ��3�Ʉ���lR�[o��H�h���0ųw�{�	B��_P "Ƅ�,%�`�,�<J���S��4P4��xI(��7��M8���:зu�2E���_�Շ%��B9�#E�#H~�k�d}��m3^"�N��"�7���v����cK���)��hI�0���u'���y�eHT�<�k�����s�@�3H;֢���JD��6X�9P�1��������Yr���T�!�ا��HP��0pX���^fg���D�o�&x���}�!�0���n:��Nni)W�4������S�w�9���2TVN۾\�>=ASU۝��$x���&(0M�4��my�8~��,��	O�(=}��8�/�5��`�����T���dh{8�#P)�.�Ϟ�>�b�60[��9%}�7^ة���f�wk�^t���o�ɭ����_xm&2�@ ���YH���T�u_*k3�c6{�"� N��9�ū�/��)L�yX]Q^��/H����)J�Q�m��d�l$4���B�o�0�����v@��X���Tl\⟝<b�|�:X� XvᛂTǡG��9�/���>J��N2QY;c��ۇF��r��մ�)H�����t���0t���Z�hYG�2�&$+���M��
�Š̑���,�zyX0�W@蔘@��
��К�j��A� � W@z�["�Z�T��ߣ=�q����{�	ч�{���{���4�7Q%*�b�IxA4�"�FF4�s�iiϊ�����rsk�}��zUL�s�IWYjV}�����$��vǰF��)��g�(�-��_��i�	-AC
�p�z�=���S�s�0ڜ�
CT�Eʞ��ѳ�8>�m�g>,!
w�X�+�ĺ,�R(H�T���K��L\\Q���U��+߾}�%1�i0f���j)�O�b/��.^vX "z��z�G��ƛ�l����ut&,����FN���@�Y_ޏK��,��KnII�Gc,�J�'U]����x����<A�x��e�篫�\��-M`���e*��D"��F@g�tttLH������`G~�y�F��L�'���^s,�������"cZ�e�ju���U%]��{��`���������:���x�h=Jg���i<I$�r�mmmh�٪�O�4گ��� ��8)ѪhI��7��Ocמ��ר5�O��uY{I�d���Sީ:Fҋ}!�EEM@o�5�9�  Y�i���J>K���S Yy�i]}��03E���^!r09�}��*\-�y-��q##�.E�F�MI���J���~�F���L6��^�aܔS�-/c?�}+�����y~���2a�qE�;�#�FU�Ⱥ��^!���?�M��F��`x]*#��K�A+9R��B�U�ooeA��\<S@%i�����.>+��h��k��Dԧ՟S�QK?{T3��2�X;g�HN��\<��^W�JSV'T�_���p��,���摁�B�!�ȏ����5�.>���qlM����#��n�_*�xSQ��p���d��W��-7Y4���~�� <Qa� m9R�xi�ie5QB=����=�t��qEQ�
�<�B o7nn�i+=�p�ǣ��{��%`U��,��ɩ�������z����99��q�̼{�i`�&�x,��%Pa9 ������)p���u��n-��w�f��Wp��o/�}� �V�,��Q!�������-RWI����q߰��p�F�%�|i�-�9����8<��o�|[q��Ϣ���*Tߓc
�}�ػjN�P)���E1̔��F���]9�E&�����O�������sO;�8��V,.�Ɵt1l��3:�K3�R����ɖۡ�7W|DAa�OV�1u��x�E_�(���f����Z�^��,��8/~
�؊�X���9�Ġ����& $�F��vAF5<ϴ������_��'_5�WiF��>l�f�R�
t���I�V��F	/ԇ!PK���E�)���^�0�����a�xL׊�[�����t۪A��[�#!~�
k*��v�������g�
����������q<Y���-t�4y�cqU����QjT���F�<���d-Z�=�Vn<�x^.��<�۷�G7���(N�q������W`^������������*�Y����Mӎnvb��K�n��\��p]&'���}�<6�w��~��b6����[��С\�)�zQr=^��i���u�)����ٓ{/[���sF�	�4��q�D�a�g�����B��h�Bo�[�����tOQM�7x�k\��?ȷ�T�r�/S�Mci���D/��O��,���TF�O��%�E=ă�h�6L���d1Ԝ����_rl�?%�G�P1�����0���|Ի.!�/���T߽���NE��rnx�L�ѓwm�*�o���G>ky��)��GK��Ѿ+��|��|h����p�BLJ���e ���b�xH~ԗT4ި�����C�a�����щ7�MD\�����Ş�3���'m��%@�dw��
�~4?;rܮ�F�R�kʊ���4��O<]�Ϲ4e�47��k+��3�{◷T�I�%�]��N Z`�Ģ��;�\�ܝ�����_'勐b�f ��Ζ���B�P�������5*2nM����Z��Ջ'�-[d�5�q�w,�w9��]5�������-�O��IU�kuH3�C�����\$9�v��t�>��oJYHL�l�"b7�N6m��G"��>�[۱ިK�w���I�,2ol�E�#���.�L�,��Z�P��&�r~�^4����T꩹O�~9E�v����hQF4	㌛�d�^����������*��Խ<[sԈ�M��n�4)c�..��{�L���h��0q�����P\+���QDQ�&��x�5�.���Y-h�� ;�m}��f5hǄŰA���R�_FV6�F����-�@������|h+h�8\���=J�q���"[b��wu�>+(�y�`jS~7������2Ʈ�b}���@iT;��ڎI���@������8�@��!?��E�lc-�����v�+�� �G��u����3����*�rrh5��Q��b�G�{FK�F ��5�=�^.4�5��v���x��p�?��يHyݷ5
���!���-i��J�Y�ᮺ�	.�X����;m�<kv��:]���`X>�i~���Fo�%���9�7����{Im�f1����پџq{�6��|��tG��X���>���e�p�w�Wm��4+�QA��F<�I��黼�u�lY#|��2�\�s4�B����CR����8�󵊟D���'���@oprr��l�������Q�F�i��uB�\��w+�S�^7+�4+T�~�UT�n-����m���zd���	�MK��*����kI���_�9;ʫK��	N�?qZJ8s�S(,���'XK\�Er�7��4p���~�ν�0����Q=��C���p����O�B���������	��l�������$Һ?�κ߳�=�dX:X?��fo��Ϫp�M'����΅Rqm?���Tg�s̟��䚴�ғ'�����3��FE�fq#O�U9�ߓfii���2�m����ѿ��t�	���#����H��߹nOD3kZ��&�4x=�������7�m��:ar�O��	��Jzq�V��.�����+�V�T���*TO.Umu'��x�k�NDZ舠auP)VfV޴�����b�tW��Ek� �m�g.��ae���B�<���;���ThƸ�:�m��K��2��~[g.k^R� ����n�̅���i�{�[�b����5kSD&qU�X]���-�X~����QY�yk���v��X�ڔXM?jŤ+�(&��L|l���.�_:yF%���f/u��ed�����i[�7`�s�$�91��}�B����Y���bA��d�4��(Ң4?��UHd��q��!=�u[��9����.AZ�i�.�
:Z��H*"kwqA �$s������<�@��%�hϹ�Ȟǖ8X�р��������tSh}�X'�1���\LVz��q/f�*������f.��v��.6�o���(ۺ|�� *6�>wZ֦�D<<�������<����"������M����b_B�(�ͽy�#A@+�����6F@$߾)����1���!L$�(q$(d�"�PV�6��h�(o�(m5Dn��p+���񝳥��n;gf��ُ�V|�GgKGg�11YO��o�ao�Zd�!%�����0���U��������ޜ��wbI�yH\�������n��dVi��>�X螃�GMJC�G]��q���s.&����b~p���@s��@M]��z�GaV}d�Y�\x���$o#��r����".kw[+o��"wX:�pW�j�L�$� �sO}�y~��օ v�=<H�`�Z�����	�\���w�j=�;�0؍R�Q6��FA8zh�5�`HU�e�m��ܪ�L��aQ:Y���ҎKr�2��ۑ�T�d�8�L#��nA���Z=����݊h�������Pf|���N(M�i�F�Wi]�g}q��Ӥ�'rΫ���Ӣ����[���C�Q����(��Nu(�|�D�$��w���S��6"���{#�fa��G�9��E� �tv�:{�H&���'��G���Q3�։���H5���Ԩ;�!m3���k��}�j{cᄅY���?<=�WٷU���5$� �m�KJ`z�=`*̸)Y����Ma����?F���G��XT
"9p�C���$�]� ٰ�ϟpb�S��%
'��7��	�_}%��'l�^^Ssk������A�xu����^;��S��'p��z��z#�W�qB���
<)uR�tø�JQ4�cwa�ɖ8m::�]�r�H��f�F�H����;��D��^��)�t&��ݲk�z.8�%�]����ؼ��~���rK��B$m�	Nf��=�)�ō��ڢ�U�~���9��G�?�h�Qn7��+٘�!֩��!fS�@�<�>���>t�&`~o�34=m���4�V� V7���Ą%�E�ʫw���fc��f�T�0*e��P��5��[��8-��"}�]�B�rt����l6 ��5�gd	�G�q_p
����=��y����(�ء�J�5>�]n��g1pc����z�<Z��i߶�Yf�F��9�.��g�Mn+�HuP������Q��~��_3�;���@F7嘑B�3��Y+'YGfv��~]��n�W�{\.lsy�y���+޴��%��)M�F;Ĝj�r3�(w�<�1�^)��w��M���k�W��}F%my�fc.�7It%�����<��3{�zz�k��Kx�ޓ�C�A��V#,�)�	�Q��Y�;��A@���J�k����EM�ՎX�r�ϒwcԘ�-�Z�@�O�zN}}���
�Fy8�ܝp<)�qqz�W)�Rʄ'��941�����=L3�j�����(�0^rv����8��,����<�Nh��:�@�><2�%|4�t������z��m%Q�75q���k������%�K�(>�i�t��6�����Z�-�I6le($�RԸlT:5`��$�y14LW3����zŊ����Jzs�!�ڭ��i�k`�4 @C�ׄ�F�q-ɼ���T������L���B'���SY�%�m��yT	_'��6v@�~2��=�f��b�j�{�_K�v�D��<�:��y�$?�A��X�6P���;S�V*�mO��u%�9;�
��K$eM �'���\�Q�Rq���8����q�[��N�R��C�^���	�er�6����씌����^љ�
SM�!�p��$�����i��g����7���su5�Lh��`�ϋNsl�`ª��*|c�rfDApˤ:O����G����':;�ٙ��qw�"+B�Er�����l`1>�D&�G?��K��ύ"f��^T��7^̳�Ч�+cm�1�����@�>��?q�u�վvsӊT30����O��c�ׯ---����i �w|��P�bb��7BP˲�佩�.�&����0@F����<,*�\*��x(s`(,�+a��{A�i��0�?#c£��feC��t�%9��� ^�U�p�����N�F����K��]�G	�Ppߘz�Pu.�=ԧ��!L�AX=��6^�b<�o��6UC0Hݣ�]7��X�M]��t��QM���^�n����[�(��n�cY����.���?���׵�BB�%CGG����ոl�JC;�S�N�+�p�ɯ�����[_U�}=���ȃ�(-(�-�"�%����AH7��0�H�Ѓ"9
�C��Đ��{/�|>��{�Aa���9k���>�И#7>j��?��.�V��=���@g��U%,����
�s�o=�l��0ඞ~Y��>'U�褨��L�:&��A&��UC����AP�ZOk�����W���g< 9`�ed�(2�2�a�;|͹�3�2kR��P�S�:X�r��Dl%`�� v��`l�&�����%���J�����rUK�I؅��y8���$n�g��<�V7Z���sO�������b�`ss�>oRhh���Ժ�q\�:���J���n�Ql���K^1�؟�V=F�+�iVr#1���ʅ.|�g:Bŗݰ�\�I+6[S)���,Ze[�@�����L��2�q�2��N��RF�?h�]��!!%����N
C
��t����j���`��� �9|i�+%��:��<�~q���̜x���]uaf�4�}��~��^�R]�~{0�E]7U�[&�cW���
�=#{�� ���S�/Ow��'���M�#��E5r��%z�m�o�7|����{J^y�}j��2";<���g!�5Ri����B�]����5�~�}�w���`�S��j�$@��5d�N\�}���u2�!���r�c.�$�M�,*��=Kj��Y��N������8�C���S�C�$�_|���|[�;�u |�~\�y5"͛&E@.kD��� ���et�qԧ���8�<�*��4��.�9-��O_n�^����꼈�'sz�T�7���(�u@�n���G&C�����GT����4�gw�(|:(�h�E�D�Z��ݨ���'��,U�+b��˵�P7a�}^��Z�Vg3�f�,K�/��>:$��0]_A 봰���3�L���q��?&ߪvb�}�%iDdd��v��v20������%�G���ڧ�{��8�$�VM2�Տ*@�p����$�kFs�cE_pl��z��ʮ�Z/q��M����n�~Lkh�_���7#���6_�L3�3���_�9Û⺖�^g�y\<�1J�ȱ�͚R���ðE��5�3O�#��	�S8�;�ni,f:T���nj���F�տ���mY�n��0�}
�EdPp�H#P?U��X1+	��Nj�o����J��!l1��G�O�^�[w-q떦 �p���C���eB ��k2|����\'�`�b��Oma7?�IS1n?��z��Z;�L	�����W�:��Z!;������N܀���g�`�y'3@&�]�Ε�|�п� [l�X���I!޵ۢ8# �q#���yPD����PR�l��A�]�g ���CCZ��)���V��b�(�ɾQ;�z��Ip�N�J27	����P�� ��ܝ�\���[�C]�>��Đ��~Q�%OѲz#]O"��]#�O��4�Ҭ����8���Xvd��9|�raŜ<@7uT��� ��IQe �"@��^^�xߗ߷���Fl�[d��Ie��k;���}4\��/#��'XR)~ݎ#����� ��K�$���glq�����)s��O�&&&���K��	�G�R����u$}�>�����G�Ć�jg/��b�Y����tjO~4��L��2�S̘������A��c���_9칠W4w���V)N��G*��af��oyj�~���� >��lDo/y��)��dʵR\�=�RNt��S\7��4(Gyf0Q�s��g����n��ٚ�(�i:���v4�qN�0�4��|&6�@L�=ܿ��%r.p䤅@�6v�l\]5�̿�3 ��?�8�չ��;X���^dw�Q�)y�o���=HF�����#|�轸h�[4�fu,��;L��FdB�^��&<�e4(�n�E��T��EJ�3y�����# ���	��w�_3�9�so�DTFXd,�}���ƆNwe�x�%�t�O2�Q���ۮ+?
��M�aDf v;x5ZeE{���=w �xxx ��5g�lp���9�aT� ��M�RQI�Ƈ�r�}����7�u�R��&���C#��)�7A�9�k8� �a㠹޲��m��4I����Su+>a�+3�kʽlɤ����JTt�Nf�0f�-Y��u�bK�a-����UD��
�;��#�Zr�Up�wD��\�D�Y��	S&��,�(U%D����p@2!z���ľ�B�C��x�/]b�֙��j���(#�r;��W�Z��@���1)��<�`�/xGE�߈`O~N�K�Dc�t�h�x�E�J�s��R@���i��n}<�5ģ���"õD�����3�����P�- ��e>�]ls�	�.�+K�5����E~�;�OX����{�%3k4g��!p��Ps�)ǶZk=�����㗤�v$?�"�Q�V�؛rz:y�I���~|��2�W�1�@I����k�"韪P1U<"��>�}߀Td��!��PתN��W�K�F5�1׈*���Pϣ	���EΨ˴�g!�z;J�;�-k��r����dU�v:2U.�ƺ����q	�?D_N�����}A�{ඉɳ�������a��A�A���6����ڟ��7�:^?�lO�T�@�S3Pǚ�|?�^i����.H���z��d�����Tw��;Q�ŖVyt�ȸ�tP��Bz�d��Dl��)b`�iw;�{Q��G�f���UM��nXj]�b�З��dk�I��Y]���X�ks��O����pǖ���7�j�m99� /�ėS��---�� [f�bn;Z%||��Ѝ�x�çCO>U.t`=���<�F�|M��ښi�ҡ�.d���?�҆��r�=�2y�2�+��L:��������Z޺ő"��!�}M��a��\i߱��8n#q�><�����$mjMu��5��]�$�1���z�ćq�~���^Z̿4~7"�����jx/N|�O7ZK��[g�s��=WRx���q�ed�Qo��ۄ[�u���x	ֽ�0PY�ٷ.bT"u+G��`���D&���j�2l|�hT#��s$����l�&��n���T��\����&���K�<������{�������5�nV�17R��A�L�|<��B�y����(Z[\��R��QJB���TRf�6h#>M��mi
v�M2;褋�ܢ��``�A�� 4t�^׻��b�_�6j��q//�-A�M�M��^a�!֪e�3��hh�1���"9J�3��,��7G�R@Gbt,�p�?x�B"�v��Fs��b����G���'����{[�a5OM��1)D���C7KLHh���Sg�T����&�5u'���E���1�����5vI8ť`KK����% \��{#����x��C1�4�����x4z���zc[�J��~dmii�u��ש���*M�[��JѸ��Eqkj�P��Ƀ��x�&nX@2"��p��(._߷�Fjw�� �}�*�3�#�S����5�[��m��ʖ�t/#dc�9u¬7�&��oqKz�X��w�Bۂ��z��� �?�D�ή\ Q��[�9e�U;��η�u�4�T7�aM��9�rU��ر��5g%P�.R�'�|��^���ѡ2��w �^�C�e3*��j�˔�S���V�U����_.�U��sN�zԑ�z�V]�S��sLT4)|Qg<��B�^�l}��y}#ڛ��mGh1��2id���;u2Bϗ.o�Tm�Ib�JJ��ڕ|J�GT�{���z����������_J�#x>08D�����;�~�n�M�$���G�k�I]�S%r��fOn��z��=-��M�s}��娗�]��=Z��#�GmuU%���Q����&]��8��I�@T�;a�i<����K^z#?.�0�S]��/���}��y#���qv���ٝ
V���Vz��då��7@V� 4Fu��)vx/  �՚��������u�%p���V?��u����.���(&��Μ��"������<���ª=Аd�=��[i�j�#/��^��ʅ��;c�@�s���%���d@=��6���S�_��nY/K@/���l�N���s+�*Y*-�l=��H`0��;b_$Ѭ(??hb�Dg&�a��r�mx�PE�7��R�
�7r1>E���LS�q\����.[���5�ky�\��3�����S�X�.�i������V�}j�������'��}S�^��K� �#*d���,���+w��̼E :ⓒ�����k1�����i��'�!��J\�q���k�5�7��:>�\����Fb'v�Vq�p_��y��\c^����閯�K4t���"��V����]F^G>����Ѵ��\�jc�8����������@d�9��V\�~��K�Iۙ;:6���+�v�d��~f�n�P��>*��F�bg��m{��o���q�S�ҳg�9X�ӽ�/\*��g*fϥw<27�G�7���!-���j��M7�^g}*�wP/A�h!
��s-�c�slʕ���1�=`����L_�tp�p�
�_���1k�X����B��&�e��'H�[��y&G T�Ҧ_� �a�ت"A��g2�mX�&o�u�n�����
yq��V�!�x�Y]�'���վ0��a���Q�ҧm�]�	�[��2P��Z"S6t���<��(��@������k����)����͒fyYG�79�� :"���%(e���j��6W�V��A�"[d���?��oj�0�Km�]tlU$ѡ �N���(�bά�;2!l�Ud�l�(���֕ ua�| 5.�� ��s�X��`S*!����������}��H��0=�13��������C���^�0�C��v	�MrLj+��@���w݉���7b&sy�Nt���6I�x�v^DB�A��]��zn���L[�����с5��7��ߊfe8�Zl����g3��O(`�V�)�$(͙7&h�$��j�W��nha`��yO����t����S_�N|N������S��z\���������{���-F�y�b;�� �����P%�4 �[��A>��n1׊�x-�5�N�m��r����Je5ӹ�H�-��.r��Ƀ9�|-UzSe'�����Н�޾=��pP���<"�Xa ���f98|�2�(�`��}¥�ձb��ҍz
(��ru��$�Tu����L��"�Nxnܮ���H���	~o����q���I�u��D�F=�"���-�:�R)h����;zU�w,���l.>C�Wk����wu�@���`�'&V��$�'� �z�4����5;�E�"G7Cͼ	?�9(o8��k�T$�aTE�I���1��7ʫ�6�}4+Zn���9��1��`�;�i^)=�׈���E=~l�Z�@�^�߅4W�:d��G�}+ڬh-��N&� =�v��%s�.��Q��(�#�a�RՁ#>�b�f�s�z�FR���F�	��d��.�)hT�A:�(�bI���W��Ρ��{(**ඬ�/ "���PB���g�U6m�'�&�9pI���r�[�zJmq
�'G��B��̹�F��OrK�W����FB�\�sT�'\�q�-7��4�?��7����c��/�9�=�����h���^+�; �bCC��c{���B�VVW�W��^��V�i�P�5������Q!b��ˠ�ܠ��12x۵'���*ȏw�׭ݤ���Xm��\KO���x���p��B]ʊFG)8[�њ��WA�w｢'�!_�,ڥ�^�V|�v(���ϯ n����-��%�/tV�s�`:E�'��Nm��W^�b��ҥ�����h5����x��|.�j�{ls�V���!S���'Ԥ�ٳ���]����'W����\�.ߗ��4��kZ?C�<�}X���MT�F<k��Yt``��8P �MLL8��S�*j��4���SC�����˕kz#���p���E �0��FT���l�����+�Ic���?�*���a�E;=8J����gAH�҃���݊ļ�(�b��ɷ��n8����P��T��B���<<�b�~(%�%��3�^R��B���3|h������X*��o�׊ �pj%%}��n����0�'��{�k��=ș��D���Bod���Q��Z��L5W|��������P�j�6�CV��'7xF0�cG&�23f�<5�c\w'�@n�3-ND����s���8��F�X��!g��Q�ŵX5M��R|8�S&#k!_II�]����0#���#b�����Ĝ���q��cH�f_I�:2agP��#[��^�9�=2n>W��j�,L�D���稰���:��VC��+Z;�O�%(����ï���{� n}�N���·Cte}�F0Ӂɵ���E�=k@hٙ��������@�`�C����I~�%bZ	�De5�ӳp��j;1�#ur`��)E ���|fR�B�¢����"D7ٛv��G�����f
� ����e�շě�wҬʥ3�h���|�����^ʥ�8�A�Ѧ��K#��.�g��������Z��w�{�����:�l~3Dc���Ԫ�����?ٳRϗ|�0>�^�f�3�^%,�6{Eo%l���5�3������O�b�Xk;;�S=��s��s���zj�Z,��z�v�"r���G�����n�wq
�C<W�B���c��u��H%3i6bHmr-�3�m�j	X�?��4}kB�M��Հ����6�\c���G(�3�A�	����`ُ�0}B��ڌ�ho�^�z@�W�׵җhO��c��g0���>t�3����=�o��ɹ�fn�iTL��ߝ�N���Jn���@ �#p���<�h���Jm'�oǮ4:�X|S���C������iy�Ў�]]mP���!OMF�t��?s����+.=���uB%����:���, 1BY����q�c*=m�M����,G�j�[d���z>-�-��]�\]�3<���񛝀���rmWE_�Z?5Po���%ʷ9�j|6��|��"��ѽ]�z�^P�/����q�x�2kTB}��!��	�H�h�=�b<�Gc'�'2�z�~0�;�0����[���Mm+e�{�u�f�U.=��+;⻟�%2�	8��+++�{~v�2@�u��QO9eU�4e���-�==�6� bv���0�����V�٣2���1`���3i��#H�!���4�Z���6�(����)�֤߽�8���8A2~��~�j�o$<����81FJ:���^"���[kT�����,�����E$hr��A����% 5nL�*$���L�,!G�V��XD:��F썍��6��IW8�Ӣ�H�AB�]�- ��&�Rg��6�0��z�s�M�z����w*.�sk7WD*��t��Qd� }����ȗ��_��H��G�+���׈��@���0��޳�<������j.6]��M_gg��.�����|�ӵ~{��/�ܖ�"*ʌ�V��E!��m���-�7�O��w�&�4܆U�p�0Z��� <�ke�>�i	�,�[��gkF�qRd��]��چw����]�_
lq��90����J�=0^�����^@l�:B���_���a�ɞY�n�Z�"�Z��3��Cm��/����C��
[3��ː���MO��M{{U�O��|3}�t�n �8c�՛�eUo0eB�t��d�NK��A��]�֤�&�1g�x�>��Z@��"�`�hgUT�����Dúz���p`xi@["$(��6i�+)q-��3���;w� Ln���+/�Y��I���{��r��H��5��C<=�Yf&��Z�ͬ�%��{4Wp/��6ƽ�������$Da��a��IBc����5�h������^/O:%R����I`�j���֜��zz�5=9����[2��l��=̔�c���l����d�}�#.�x[`���>P�Ga�l_�#S ����9�
��G�{�*��`E���x�^լgO �	��������nb�Զ��Fм
�f���dԫ�	��Y��"��G�Ɋz���$�Dtj�w�uw�k%�� 3:d���Vy6]�f$�/���o�J$%� )S9��}1((��i�$��߯�t��=�2�XGG^ri;M߬O����[n��a�LTe||�`��zQ���(�S@)� �4��v��Z�u�����'�ydJ���4I��I���1�>{(T���H����q��x��Un_���Mne	�M�k@A��8E�/I�~x�C}>{�,�m��"�X���B<�29(�>@N~~<2y�o��^{e�(||`o_���K�ug?�oT����oHO�	� ��D���iNe�c�`��vuբN�����z��nKG��#M�Բ7"�|�.���t��]g��3؞5�
E��|!#	���ۼS����_s�@r/V&���ܰM����p�u���#+7�՞�(X�`[�㜉�	@�f��!v���q䌺������ވs�=�l�<��5}��Z���'^��6l@�ӏ�ٰk�HX��TT+�x&��Qw����RS���2w�b?�d*�.Հ�Cl��-Y2�{36(��Mzz�?5ï�u$O�[o#� ��� 7Y$z�:6��5P��i��5J
�>���%�
�9I�y�bk �}RNh�G��l4��:��R��e��C/���Pq_p�����i?�����Yu�
T)r9�zl���� נ��������biY�#�UX��R붇���A���D���3򦍒���@���I��X���-+Fߋ2m�/I�U�=��	� ����	���?�r"Nkg�0�Y���l�qR�<�{�%�&oU�f72���Δj�*��* �^8�+����}'e��R<ڮH�ۻ�c��Ѕ��l�ł���o�īh�Ǖ�h���Aq��_�4���r���X�;G�\�v�X+�n�}�$��84
vY��1&X{�t�@�R�!�����~QvK��-����h
�=���C���@K��FPJ�<���BZ׮��_��O��Yԓ�k��c����n֌:4=��hd�O���V<$�äTop{�G���]њ���rp	�������I1���VO���(��bˇ����9�N>�#�k,�w3�6�>&^��p��,�3X��@�;-.m�A��DȚ�$�V��.��PŲkW\��W~�A�庠r�*Q�u��f��Ml�ºE���IV�ʈ�̑Vj���0�3���!��l;S'�ZMS�R���j�OfhV'#���<��}�\�l��m���oC�l�����r�D����+��-%���u�o�~�ݨ���~�Km��ş���=+���>�S�7�b��7��������Nt�[�<�ǵ'�+��/<����P����A�2�X���ȹ����V���?��6��,2�U���r@{"�v��/f����#ã�Y vfZ0�#ER��f��`�qk�<���Kq�� �
^��mju�������׿W�VYw�\�e���Q"�o��E���N��4\�Wt���9e>��&�_�I�N��m��V�wz��7ʓ�w<�g��;q����,�IE84�=ux�I=�����Q���8��|Fl��@�Mg5RH(`�Qe|ʶ����1}�'������C�� sKq���)Ɛ�м9���Hبk�ޭ+���2��;��!�@�m���X�)7�X+��#ރ�T+��-���an}��z:�������ig4���VQC/૩
��+��/��Rq`�O�,k
��6��[�OYk�i�d�e#���ꞻ�͒���&�Z�"p-���!̫�l���&��ZM'� $d$���D�N����w�".8q�Q���
��R2�G�!<#�E�A'"+��ǐ��N�٨��%��L�L��f3A�_��NO��?50�/ӑʢ�lm;��LT��]�̷�5�v�Jس�N��Rc,>*B�=��|ʀ�R�/�-,��j�uZnZ_/�J��`_8l󏊻k�Cu�O��UOJ
��H��j��]�����e>k?
Kih��"Ǵ8���ɅV5�i����o��{��n�>��O*��HР R��BS0�������!���߳ ��)������c���C��-���}�鞵�ؐV
�1H?W�䁶L���i��g����0!���!#ǲ6]dJ���z�n�������٣�$O�Alc{��P���f��vG�����uš����d#�P�
5m�w��h���n�U]���a���k��~�3���Z�N�_���=bE�z����x�WO�8/�� ��l]t�@[ ���T��3Kٯ��.S��<e�������JD�x�������48�uO;��!�?K�{��wn~����PMٓ��*�\��Xx�vR$�kYw��x�J�w�&{w�Dw�(+O�A����>�m��;��q1�j�(��{��B�����(���u�b��Fkc��<�Vhj�P%�z�[/���A���ԋ��!�cLw?׉S,0�6o[8�����n͒<�� �~�.*�?`�q	 +(!�����������>ņ"sg�?e��N-�/��<��}�[^��F�P�3��Tz�T����٠���7"�w�N���ӻvǵ'�i#�GJ�H	���_̳����V;���R��^#��4�0��Y�H�b�vv9GohU�?�7Ɛ;��Ɗ�F��N5��ߨ�sP�/j� �ķa����N4W*��X8t�ޱ�x>�I���m-��	Q�J�={F��i? \��Hrb8p���e���P���`K�� k�[� � o ��[� �g��@aG�^�=OΗ6�&�9V�̼(��/Xb��_�D�:���ݳ��B�hu��{��~>ɷ��2�}e*l�W. h<��/@��4�Q���ރ�耂t�j*�n�L+����n�>y�\�W�j���Pzd�cnsC|�>���:���-���p��'҆`��鷏���_�C;Ya����O,���^ �Wff��Y\��D�PSYlHn��V�C"��A���ډg��:-���:���9�k�ٞ��oj*�k9�	D`K��N=����+�����x��x�:������4$.�iL��_��/&Y�U����S�����F�+������t��6����m)����1��>;�,0�UXRRK"���Y�3y��Φ*��È'�q?ל}�%a���,�}�=]-���YV��D�q�)/� �<
�|:&z ++�Vo��<ǣ�-�p~�����捍O����5�W��i��C͟�X��~��赔T�i�N���s��ϟ��b���䖿'b���'p�@A�.;���:���m,@AS6_�/XY^V�8������ox��o����*+G����Y�C����Fs4��߫�O���{|� ��"�zN8j�#�{�P�����j�}�F����	

�ON��F���,������e��͠<c�a�;+�!��_�� ��௷��L�������\��*+�Am)���{�/�'���If檪�����<�H�spp���w07����5���J4�k��F�YY�v��������������:��NVCqaaH�إ9j���(���Ç��]w0hOmy�����ݯ}����H�,//�.�GB|���e��!|���sT��Q 	�	�����L���3���N����   ����h�hKuh�!~@-�"��\ o	�엿�P�;6V��f@EG�FA(�m��es���('�XCK+$��,p�\�AAA�#kDw���^P��X�&gUK$�SQ\A�����ܯÅ���hmƲ�0��?��r�`[W�8gp��37���C7跞)p�����U�����>���γ\{�H޸[Q��v'��oj����o=��wS��&�������=�n-ߔr���"K�~�bٟO�L����;�s�����W+�@X<�i#��9�P?1�N�cP8�*���6��n�� ��/�q[�l�b�_�]�����<�����54���~����,nթV��X�s[Z�V�+aj��T�<W�S��hv�%���Y.�'P��������L{�m��8ׄ��yDm�/9�\��R6a�E­ixh"��5}k�̰sWcB����f���ס	[�t�Ԥ�%7$�4���4E~���9\�"-L�K�h5u �j��9`�F7&��3|���0��v�ױ��Nv��cw-�����q�I��~Rҕ��I�Q8��v{��_^	��x�BR��{��L�$����8+�����0�u��e%��`�Rp����zn�n�@E��eG)1m�������i\�#��(��6��@q�ݥ��;��R�O�Ȩ�l4E	�ye�]4��1V��Ox��E���m��2y�(	S��FS�� ��-v���,�z�ܠ�H��_$��)� p˅�o�����w����	������b��)"	��E��F).!b�y�]��O�u�=�#>G�);�S��5��:�I��c7d��m���_��η4&{h0���w#B��:l����K��<<<��� }�4srr�z\
�ܘ�:8Jp�LBId-l߭�o��>4��\?��K�$y�����8���P����j��t2~�NG>�Q�"��<�����Ԫ����G>�g ����LjFݳ�f�xC
g:Q���1{@�)Y� ��6��,����Ҭ�x	�h�C?lg�7j
�TNE��8M�9���ic>Z%iT�D}O��J	�9��ތ�]����t%�۷^��K@kxt%�>�
^*���2:
��� �PmD
����|^��b'���se�eR���'�Q������0��Y7��]<He�ڶ��%K�L�T��۟9��ok?	.(ѯ��_x_9���h�a~��-/�V�mޱf`���9���Ƥ�xp��@#-���k���4�Ż�ѿSU��!���R�נQ&լ��\�Y���[���b���{���������+/K˧�ۋ�@� ~�{���3� U.ܭ7�qY��e�M��}���#�����Pb���/��պ��5�4=3<�1�^��E�ZyTKD��Y��k�~E���8Vk�\�dg������
�;GR�"�:���`Q�{��*�v+�w�L�N�����DWJ�4iۭ��j�J�)�1��0�j᧥����~z+��N���KD&rЃs/������R�j1�N�{s��K)>8�Z�g�������q�J'�W!�KB����/��UXN>V<����ɸq��P;�:%I9%�i�˪̓0�����r�G�F���7{5Ggt��n��jH�|{�}O������ ��g7k���4TUo&��^p���U���w�����D������3f�S�)���/�������k�B�;����f�<�=����0�y�3���w*�{�vZ%��������>�\��V?+{��5��򇲘��jhzl-�������2�d{�s����y�uޣ��|���'��q���,Ͱ�f��j-�Ct+�RˢU�����a�Oz�$<���R�ec�9x��0偬c S��e��{_�R�?Yb����I��3�I<=Z�n`Ps*����] #���(��u>��E��zS�{��k�����NSLq�텛�_=��zs����w{��-!!q�8����dk��'��|ƶ�f�e]�b+���)�H���:���է�S=""wF�����[߶��?T��j�4�Y��u%f�o�K�^������<��t��q��[���!S�E�J�\�Ͽ�����/�����n���#�R�ae��fV�BEK+H��ԝ����������0;���['���^%B�ʌ�G���>�j�ϊȬL�ACW����n�wE]��t�nѲq�y���/ɕ�"���wŗkh��EЉ|N	�egUp����@�>�ק�>�����w�Q�8��.wETݵ�]-p(3ߎ�t�?�x����%1�ؽ��;,Ȧ�x��f���u���}+���t�9���o�]�JW����ۙY���tt.(��JQ	a"��Gl�%�a��Y�������+ (�Ɗ��T�]��R�C?�9���|�]�Ue���nz����k�Z�9�S"8`�-�8�%�Y�z�����y�B|f{�M����[�M�{Y�y��9��W�e����h�sAfJ��U�Ϻj���D2�}�޽�A&h_�	
���޽{���VQ'��ic�F���_f�э����O��e;��^��#�Qq�9�)*�V�����C��,�����c3^P�/�
׸跻��dO�Д�u���/ɤ�ۚc�=�6U���5ut����U�H̕D!�ּ5b3ۥf��4i���y��k�ќǜK4�7�`�E����P��mP��fpT%�������	qu#[d^������ <�� ���c���!�xz�������:}���~�ue�y�B�c�h�o��
�g�������r:x���ZvN�7�s�E�()�
���b�����s	������[a�"$O�kT,y���{d1W)�)�Ho�d5ɉ�5���8�ZtZ��mf��[|�w�Ia`�"��;ˮ��'R�m����'�7'������6/�����-�e>���O������P�- 
�jrʿ��^K*:A[cQJʼ��D��2.�JU6�M]QJ5eQ�#-Q�e�Dԉ�e�.o5���;r5�!������W�o.���5\���7���y��$��^dq����ʿ/����*$�ɕ4��ҷ`uu�)��m� ��'���+@���.�+d���DO �	]Ee�*�Yi��G�������i!��r��ȝ]O�Ŝ�����Uei�a�a_��D���d��4d�^a?A�#h�b�$$�]XR"}�i��r��ůA�2S�[oO�������Cg��qF�b��
{��m��:2Sζ�ʻW�V|7���{T���ߺ9S]�#L!�9��-^�*S{�>��j�#����0B���Ĵ�=RW�z�����O������dɾ�������O���,'�f`�g��m�U����{i�����\�x����EB�)���9�Ⱥڋ0�w֯���3�Ĳ\�c�f]f���	�OGy�<���Gh�<R�|��_�ȋ��,���47�ĳ D�@�m�{�}����-�C��ؔeZ��a�'6���ڒ����|Y�x��
Ӭ�| g�"s��j�8�������8O�L��ޕ�������i���iH��8�o��E:��W�#�Yd��&��=ʵ�{�15�I������������ª�5��SM����ݻL�-E�� -�{(y5s��%��zC��y��3����b�Ɠ�V�ד/�k���M�Dڴ�i�ǚ!u�WDu��u	�察
��i�t�����ۻJ��(.��=��
��o�H�(R!7KlR��4�p��t{�ɞ���[ݍ�<�Pվ_��em�f����6"�XD~>��k�9@��prp<24d<"|%�BIy�K��
g�I��~B��`��\���~�eE�U<Պ6����3ۯ�c�'t,V�o˒�|��B�~�v/f@��^�1t�rD�����\ĸIx3Q�����e��?~J�'è.ob�r���kʗ�\��Mk�x�b�@��}�G?L���11ީ�z.��MK��S�`���7��k��K?Wz,-�lnA\;Q�:��O�ͺ������IaJ�;!B��׏~=�m��9�r�p!%(��Af�G�Ї�&�W�'���K>�+ڟ�zPJ&��x��溛�#�Ȳh[E�[]��[�7�i�TxIik���[Vk��$�e�A���Q����̣�o�-]�=蚎f�/�W��~��={4�y0by��(5�ğ{?����}�I(��}�_KfY��0����5�
B^ ��c~>IJ���CH����NM���MY7�yۉx�cj��̄A}�Q�_������!�xJk;�u���%I�R���lH#���D�Y�K]8��f��C�|�9��W��e�v�6����9`L�X��L��h������b �]�	R}��o�6z����U��R���Ϻ���yz�"pv	�H�ߠ�485�ٯ��敤��8xxd��%�^�
��#'�[a/��Ǵj&}y�lS;��L.b��0���sJ�l��FImMO���vI�>0�:G _��-%}�G����'mY)G�9.��;��hM�Ic%��&
T�P��m<5��V�D��d�M�+�
��~"�c����{|�w��,-�Î��[]o)Z����)ۇ�$�<��C{���y�,n�� �R���-��*P��/��ԥl�}���^��տ뤪w�����y�m���W� ��v���j�V�����{!�jg��p�2EE�o%zu�2�
�ߖ��й�"�5���3���ƜI��Y��
j��ݷ�|�N�o�U� ��1�p_;] �������L3��S�Y�)){�m�U�B���1���ju���V�)���?;8���~Z�٠���\@ ��d�����܏��.`�ZV��x���\��_:��k�����jh
�����CoH�Ժ����uh(Y'�pc�顡L/!J�)���5v�����cY"�[�4IS��%�^)��6��3PL��ͼ+ۢ��xP��?��׵���z�1�C0wA��lf":����Đ`��9�QW����S�R��e��9��ش�"�L]P��4�-u��\w�#� L�2��T��$�k}��X���i�Q��9�x�����/�g�-/��wtv>�b�I�#�FcD��B���דfwf��vQa�NS���"������c�=��-�f�
��bX��� 5XP3�	S������w�Λt1U��M6{��NtHH���d�z��8(N]����/p��Z-�.?̇\kT��2,s%#0�i���z���l����N��u�+W(]�ZV羸U'���1S�w��R����xa��]�ОX9b�(L	xz�3-�Z�:���=��u��3v�E�P�^i�|t˥g��>��K_�8>����#����=]|���\��36#������9�����;N�O��X'��,���c��&Ů�	#_�(��;~�A���p�Ж5}���~��1	t<����2!���V��%X%Z�bm�GlIn���b�����ȳ�?N�X�-��k��Sqñ�ۤ����*��:٤�b�Μ%��g�!���B��9o��Q��lR�I����v&����#�0�������΢ϋT��(
����]�'���W�c��� #s3���gq�7�uq�(����wUM�=��'�E��`)���������긨���A�CJ�F%��TJ��;��2�P:F��C���;������?8�}�^뉵�>���\r�z9�g���f���0������,�KU1M�X{^|�k\������~�AL;dTHgb�����/�-1�N+�~�D���R�F��xK�};��ײ�ʰ-3$<��NL�rz~~U4��_3�Kwމ��}~RC���7�w� ��?����k|,�E���	TR��pf��r �K�}EF��wQ-*���F)��lug��K�܍�Yat�
�8�LL��]>�� ���G,�x���߂�Z@�<�4�9��W���]����8�Q��0��I�����U�h�z�؉7`����\=N����M�5Ȳ�]rh��d���PYT]8q qp�:u"���>��N���}3b�|�S����u'giG�&I��Z��}ȵ\��b������C�:���r�����6s�؁'Y�bA�i �6	�Z��W��<���fo.;L89�ޗg�?�yS�b"O�0����'^[WWn�E���j�EB�F�����	~rjhxE �s*rb��2�$k|.��{����b@ԙ�r���ҧ}��`�i��xG�&��#_Q�x������|�B<��Lg՟�Z�����	��8����(����M�)��!�Q��ch�z��:7M�ýp3j<���x��T�����W���+7���j"��f�W��m�W�\7��m7t�����w��Q�k�$�v�7��xY�HA�tW�˨Ev��HCu�[!���#���!��~�+��eE���W�=�j���Q՘+<�9v��9�� $?�N�v)����$���A�����ŷ�&�jq���N�s�^���t�Ղ�z`u�Rp��?�=��S��qU!��{Sj��e�V�k�A�j����#{`��_7�r�هA��ά�l�x&R�7 Х��U���H�pOC����X��t�E��ן_�����F�Z���/���yыɟ�3E�=�����g��������D���rȍ�N�p�}+�3�@�qNif�Ә��k����*��v�"�#�d�!À�+k��@9%��¢����G��� �nǎ��K�%]OҒhܰ]v�ClLI��9�UǪNPd*�!�	f`xo����)��j�ow)�}�0Z������������`�G�DZ_|&���69�`ܖ�c���oԏ����׮� x�ʤ`�����@A��ϱ54�����R��%G#��­�S�FE�A�����'J���b-�a8ڸ����Y@Ff�)ī�{4�.y��|��"iŹR�c��Jm覈�N���ؒ��s W����I9NH�e���=��SW�r`s��?�$�'�Irer.�,��_����IiiQ���ii�i?�p�l�������X���W��!X%o��D��["e2�	e*$��K���w��G��I��e�t��z	BV� -�j[��#*�$��uZ_����0���ݕ�gë5R8�(�UL��j�(�?�I�9�Su?uf_�@6(LT}�����E��op��b�e`���2��q�E�ޱE<@M�5����� �k�|?@��8���<J��ȁI"���D6g`����\&}�W^1���X�&�Wy?��j��I�z��H�����9�T|�y�y<�wVd����Mp�dT��=�!f߬똨
j׈����]������[n�G9�ͣJm�lr@��A)a0�e�Nu��H@���LV����/F)N
�
����բ�8��׾:$��!E,�����Jז�ƺIݯH�����閄�I}�⦷ �t%]���n�dj�%�&���=!�n^9Zʉ���P&��g}�|-K�[�@��+��I�=?l�V�1(g����c`/1�L��󽘰�w�"��WM��1���[DkJ%�$��g
a/P�6�do����b�u�>5�a��*����~T��a�ogs�y�ʖӤ\�@JN�t㐂v�+��ʤ�h���A`�[4�9�M���đY��]�!)����P֠��aϱ�T�4��G��U "���~z�_�`j��@m=����]z��c��;��ǂ�n������)���hh�72��Ѕ< Eы�	�4�{	i��x��$��+����V��*r��K߾�-�'#9�Ÿ�?	������H4����DQ�5���mf5�~�tݶ'n�XiF��N�6�����lR�)I[Z��]���������!*���~W@i�@ �]Pڇ)�'I-�1:Óh��WEK�.i�WZI�>#?�!�"7#x�
l5U?�J�i빬j��2X�{ȟ	���i�N��>���T�a�@
��֓��1��C�T�ꈦ��nZ�y��p�Wt�����C�:�YYh��x���X��$h�d&{�Nqw
�RtZn�|��Mv�UvC�n�"��H�'y��������@S�uJ&�N�[-t_�x"���"S�.U(�݂?-���W)�mn�����������k��s��N������44�`��Gb�L
(M���I�u�'����7�����cn��fD�zVM�"1q�[d��9*�o�dA}T����B������p�nu
�d�*λ�ºո�M��1X�����!��A?���W�kb�&�``Jɝ�M�ZO2Y��'����[j��]���>]�m?Lz.��&N�*j����Un?+�]�Y�BD��?���O��X�u����2�ֵ3ړ����}��ʔ<�����`P��q�q?M���)"�G>���9�}��$L����(��Rz������7?Yp��cp��C��`�J�`'*K��&|���|9�Wd���ٽ��{���]�C܊�Q(�e�ζ'�M~0������:ܐ7��IL^^�\S�����8�Z�Q��F}����i)�p��qkLfe{�g!��sf�tA�D#�g�z<��#���b�u�6�4��%%����� '�c�ꍠa�}�@{��^�D1G,��H0��a(	�Ltr!�s�z��*��"$�c8��I�'&<�H���iC�iC�������f��g��j��\l-��YiC_l�=P�FSt�P��f���	��f�!�\o�����ˑ�p���B�w����bl&��VT���\6�\�����_3O6(ZM���K~��+-�P�C��g�|itK���^��z���Mw0ڼ4��O]�O����Ǔ��� |�Њ��E�I+���9�����eZ�W�­���V��琏�T3tќP2�Z�;o?�����5�D|��̀��#��Z�\�pp�0�"`�H@����RP�������W�����e �jz�$��!Dt��X��e������������>��:n. =Yax��� �����n~�P7=,����p̄oU����� �?�#v�?����x�S�K��ǌ�O���{�P���W��|哺&VO��:{"�s5i_��^8����s}�H)i�p��1��Ƅ���n�1��^��������ff�O��%�� Ҙ_��)���V���Mzv.�Yh��,���}j	
�Nͼ$��)��^�qM�Ɯq��<��-���*>HbV
�^A���잻�D�b)�I�8�! i�X������s�,��h��}ʸ:��`�b��W�n��>`�λ�x�8F}0ܫ��Gy[Y��Fs9y�-6�d��@��t7I"lDB�0k�
���E�Y��;[�&�3�m���/�0������=LǱ󢹚S
O��C�'UE<َe>��F���UVr� !��t��wT�l�-�X�1��sd��Ao�MG�X!��r;��le�&�3]����-��&:9c�jD���Yfi�U��B�r�%����o��K���^Hym/࿖��� 5yZ����L<�Mt�h:f�xh�U����>�ӣ��]���Gz2����8���;T:�j>����Z��ޫ���

n8�gffTc�g�M r�9`j�/5�*�;g��,�^������%�n��#ב���Yg�4�f�]���\@��}������w����F��9d��ĉ
q�����B��ɤ6/2O�@:�U?���I�4in}��0P^�S�����/��/��G��Y��+��~��ZΥN�A�X�Q�˦��]*@�s�o-��וNYqd�sAE~Rh6��i͚�HO6z=K��p�d����v�(�US���2qܷ����Mw�a��O��g��j �/p�4H�7��d�Q���r�l��Zo�_�'��v3� ��m�@�4x�"b����j��<6qr"r��~�U��PGZ8[�N��4a��P �� �Y�#�� �n�֮��Zg�����|>�~��q�7z2�d(��EĆ�+c�{�ړ5=�'�Q�9�3I�w����-Tb�=!�x��ĸ����s��w��-hmܤԇO�~a�Ff�&6-�D�(��"�t�m�wc/�2jj���^6���y�G�dq�po�+
 j~�q��T6F�=�(āÞ�!�g8�O6����I��c��_�0�L�Lz�X�˲J�[�e���2\M���aք����Өyt6�6�Ǥ�[i��c8�j�(0��x�@~6�M�2�}Q����hJ�ƺA�xĊU����@l�θ1���g_sG�UMaPq��s��v�S��G� +�]�/o�6w-��/�l�|߲?CJ�4�}w*����n�C=Oy����eZ]_0呐�;c�Vz!d	B��Xfn���3RyY� ؗ��a�/��{֜�fu�%�F,���Ђl�I���;3��	��~��������М$0���W�Y@�sB���rcst)}X���W0�����s,ʯ�䤄��# 8�
�����췳�J^�7�2X���!V��Y�mͶ�v���X;: Y�����a�떵P>����<{{��e:"ޯ�'~�
�	I��K����zڳ+T[<]y��r�G�5���D^:F�t�40	�0k���'WK.���)��;L_�J��=K`Qz �J��ڃ��
����xA5��r�Skv1�����bԇ?�v��IW̄�*eq�����tw�b}Y��S�o �_���]?��}g���@H����{��A`B�	�}�S���L�K���
�"�����{�����R=Yr����ԡWoP)�Q����/�Z��.�ݲx���HB�%
�@��؍%E��ӄͷ�.Jc �����X�|�vy���w�r�a��c8����y�&~/��l�7u'�S]*�%_���MrK���p�r�zLe&z�Dׯ'���Y��=.))���j錦6��A�� $	8��;�!`����=��v�`}j��J�|��q_Dla�r����s��P�Px�ڸ��#�s�e�:�{%#�	y
�mnd��GYD�Dhm_{ٞ�9���<0k�J��M�)j�M��`�\�����e��HA}�'
��ĺ�2xhN4W=���C�H��@�����Ty?,o=-�h�����+�vY�����-�8���ҊT
���Y��G�����Dj�/����?��őI\�g����?���&���ؗ���X�/�vP��u2����*�;&�xx#�� ��c�S,i�R���-�o^�n[CY% U�S����WYm�=o5��
���-�Ơ�B���3<ե��ԝr�Hf���������*n��M�1nv�*c�K_ˌ`�~jީ�#Eޡ�4�ƽy�����t�C̥�c���5�L��z�C�;l�7v)�n��&�վ�_�w� ��(O�0P��P�h@�0B�o#��*9-8��1�F��
��l�ʘ�5m��un��Fϯ� �,��K� ~l�C��[�?[VxL��n��q/,����x���~���!��4����aW�:�Ô�v�����X�� `a���-*��Uo�? 4H��Tr~m�h��v&>ea�b�-��3�fF�F����Z�XV�2O�F�Q����,<> L��	�o@�&�'/��6��S��a��Ao�>��6O���oH��І�W��o:β�x:>��Q�>�
d�4�d�!$6'����䏌�G+��K�h�?\}Ǘ�i���PU�H.۵�����>;/z,�|�	�V#
��=��M��a(B�q?u��((��Z>ʫ����/�3?%��,+{�T��9�1�q�.@��{aa�����@�2�"��uCY_Ai@j�������=��z�!<��4l#/T$��}�^�k�ͣ:W.ÇJjo?G��b�=Z�>���/=nWv>(�p�e��R"�#��O��\i�E��*d���5M�q~��0�����o��̪}O����MTQ�w�t�L2ϛ���Ƴ�]DٲR��H*u�U���D�Kl��P'���+���鎔L�N2 ��Q�_���I��%~�=��L3���--4��9���GAA0�?O ����t5�k;��G�qTK��^�k����b>Sܥ� ���2s�e_��Gw[qrr��oO9��I|6���P#��B��!���{cc��h��"��o�^L�!�1�x�6��P�r-�nʭ��/�^Rs��`0��.=8@빴((�~\��IVE�\�ͳ�/���eƸ�^<�n*3��ڏ/
޹64H���d#�"Sw���w��p}`=�^v4c��/lohWRP2E��W`�T^�c��D�?�`�.���]�=�g��48f�����S༂td*�|;�!�s�ykp���M���=�[��"F)�l����"��8�@��*�i�u67��5�t�.�}���8$DK���#kv1�	b����GKB��~�mg���&��A��csF~*	@,cOj���L �?��Tʡa�+Vz(h���o����r���Aj�����>��M����R�_��^E͑[Jy!N	*;Jd���	�`+� ������3�_�w��ޑ��eH���hc�� 	���Gi9�&b���WN/�j}��Z�����SJJd��u��#��ih�/
�5���o�\s�)��]��7O�Qx�l�>��{�>y��hn�@��؂��?����w!N�~+��F	0��d��<Q~x��n/�  �Il��
'�6,t#���O��HQiF��yA���p����T��SC�����P1�M3��cG���V2�q����/�w�FffzQ�:��ӭ1�x���[IJL���H��A�ݠ�̴�Pt��x)�x�9���E;�_�����#ޑ�^�; �$�!� ]�f�1����{nM�♊�#pQ�P�Z�3�o�Ҕɘu'�a��[�X�B�qǟ���v�~��B�T#��E=E�i�:��� �/`�|_�#���6�>�����(1_c�F 6���2c��vؼ`nnO�p��&��r��\X!`�޾���C�hϠ� �\���l�^�GIt�|.66p�;�x+鳕�:V��ĕj�	�b���9o����ﰠ��޸
0/�k���U�0Y%粦m��dT��Q���N>��;�J�ME�+�}���ո�S�/ՂJI�h{�������t�����J�x��G؆On�����ҟ��\Y�}���/��NvZY���cTv!GrJ���|tY�5.E$F|��)q��{���o�p$�C��	��Ce��̻W�;t)���D��1��ґ:>߄W̖����٭��I^��U���!�_����D�d��.�]U��Za�5� ���H�l4Тk� ��/���4N�tA����U^G�h���D�_�T��,��(��;�3��O�1�"Re��H�nn�����a��:�TY������=�_��z0��YT~C��<�8~OFN�w?�s�� ��}.�b_��]�hǃ����5��ZD<��!�l���WUx+�t�Hp��D�̌[�#<��L�5�����>X��WJ.d<�[� ?���TÆ4Ṃ3f��^؅}�B��F�t�[o�ܾ��:aQ�)>Ⱦ̜�Nyſ/4�A��q4g��,f�P�ł�# IL˿�.�<33��w�hKۅ�/�(HJ�l���$��͇�8o/:���S4�`'*}�sWlY�!!�����o*�z΄IO
��-L�U���kBQ���Rۦ�� %U\��U�������J����q�_�����A��0��"���tdc_�=	5l�	<��Pa�h���Ât�b8��>�/�2z���9XM����e����Q���v��M���L.d�@=����4`�⮮}iG/E�5����-S�/�� ��h��W�v���H�\ �)a_�9�7<W4
83���;:�]���P޿A� f��ޙ���`N�瀩�lo� �����[�lPb��$���-�����!qbbZ$�ߔ �{�v�,I��#& ��#e��d .��]m���FȄ����z������/1�G
@d4��3 �(�D5}wq�SE����PJ`DG}� ܼAl�`G��/����!Nv��pynv~��ذ�}���gn�Sl2?-oO�YAgO��PP��c�z1��Y���N��A�~˯C_���&�?=1rh?��"�H����]���v�FOM�L�\���_�~5o��E��=����̢�!��My4 P��ֱ�$��3݈�B��"��O6�<jڧ;0ѣLv���9�qC����+ki��I,U�~�ϡ�6U�ܗ5����Exݵ���V��]?U0J@5��d��;J=��:���k/��M�<`?*Cd�,�k�$0z>�b�D��]*k⽃�" d8)�!���!�C5X��<'V�����n�,��f�BQ���0�~�����H���=uAzJвnXzŴ|�c��p*�)>�_��.׾�Che�r�v���Tl�kx�<� ��f�s/�Ũ�3C�ݾ��ւE�+gt8{A�R�h�*It(i���$�1}��xm@ʇ����V,����>�.@eL"O\���F�s�8!>��ϜzDѲG�Ee �T�S�������^���wo�d���=?DF�})i=����J�y��N{�������u�_������V؝#�iC*���B���Kvq������.lǨ/x�_7@Vg�j��tP��s��p�/_����M��О�܍G�K���1��ė
��5�� �J�'Z���?ܽ�4�׽G�lx���A%)ˏ��U��H�9���W�G�.rh���9��>�9�� 8�ǡ���b�Ε�D���c[
Hvܛ�.��%�U�����{<^:o0�����y1�����W��	�>����ͼ���6�-l��5����;6��6�U�D@7r�X4�ڪi��M�
CV ����?s�ܖZ�qFܻ���d���`#�(��Ξ^Y �~�#�@�q�#��X*R�AǞ1�D�^Ķα�eP���@�cf&�Q�D���.V��`�;�E������'~�b��ܗm�����'�o�^��I��yx�*���Ȕ���=�ѳ�}����Q'����j۳gP&��\�,?TC���V�RL���+@�d���-�\�_u��T���*S�w�6�it���Y�~d�^�?g�5����}��o�ɼ�p^�rm������;P�f| ��0���i�D���qr�m|���?�1�;	ĻRMÙ��3���XU�s���J�������Q�ß���ˡΨ�1��H�����1�5��a�jN��F)���7�,5GJD�k�d����
  �a�t��V��.��CS�zrb��X�~d[�3
 .��<T�(

#J�jL���ۨ�ԕ�04��G��w� سl�qzIS�w�٠�r�S���	��M�
}������R�{3�hf��[:���������h�^��������0B��̒7]�}Z�bM-�K���l�9�#��G�O�%�Mm��]�_$n��1��.���:f����:kj>���{U��\�vmg�I�U�ؑZ���ğ�<�6 ��k���DOk�#(�;F�] 	�:����Z�9kK(��c3-��|@��5=��i�Wm]� p�V:�?�?�����f�G~>6�E��]e6����B\�)���b��\�Q��k���t��X�k��'�	��� n��&�&~2u(O�+9���&�qQ�����g�kJ~|�s
��2�VLf�ש�֒�ƥ�����Y�?S��B��G���F-#��X;��~7O�T�7�d)�����[���o��C���
!ɱXv�љ�!I�J�a�񵄀�L�Э�;&�	�"Jw�g\���b������I�ܴ���vX��Kg�&U�̇,�{Q�lN�Ԍ�X��{�=�kx8O4�d�/$%Z}���4�a+���]���|@:D��<� e������z���:�2�=!��S�co��|&SO�+�
����XUmrhSu�����.A�6FDhA�A���"e1�OgwZ_"
�3p�\d��|�_�/�8*��_���J݋�2K�%{a���8��v�u�[��`&�/E����\���;u`�e�r(�\�-�(����op�l�{x˪���O��q�,�����x�*[���_��������C�:��()P�^����~�h �>	
��C*�)k,��Z8�l+C����ijIk���k�=@��K�ay�C =P�=nX��2vc����,��@X&u^j�r����"���G�x=���>F�,s�&�����RAC��U�Y����B�%�{��P�D�q#X��g��SN=����u��8q������������y�\Ũ�W�e��U��'��o	@�ii�:���xD:k��[	�<�#��}h�Wx+�-�=?�v�L����(���3�� �hI`��D���?s�F�u������k���{ܔRa���$,�t�}�K�k���ʱ�$A@�V��D��� ����q�.�|jJs-}�����M�K狡���2uO�ߓl�FT) �Qr�6�\��v��� f�C���!���˩%�0��`rKd�I�;���e�����)�,�u#k�q6���w.ϸ(�dp�wR<�v�s� X"���#��Г��� �4�HR?$�[HH
ֲ�*��o.,*I�eV6KO��t��.���ELdU{@�2�i�.$�ԝ��B���t�����=��˨}Vz&u�1�J�Kª~��w8<�E� ���w����E5
1-��E,�bt�OY���۴�lAV`L1�G��X�֏{c��P}�5�hՊXOZ_s��Kql��
�5`s4�9��&���_�j����)��ȃ:�Y�꽪��R� G��G���L��'���Ş]��=N�:�}~�%g��%9=҅�96.s.�E��8��i�E�[�Z����?���7�5���g	c كȡ� ��䀿;�%�S��gR��y;��!��WOY��:�7����\o+NY�����LU���ݫ�_�&���[���c���������N6��TY`�3����
HL8���P��{t,�-��w�-�/����~~N�YO�T�j},eϹ�s��,̋�]�}��7���;���]���P�m�s'H�{#�����1�?bEz�xCrp�ܰ�d=~D�qc�UW��=*�*�s5��/T����m\�x?C��/�a�f���d;��N �x����.	u�n &�DIm�wCɪ�F߸("M�r����~��!�����:��
G-D1�I�r�4�xJ�OH�2�Q�b��ț��[��=q�
$@��^�' av�o��L�+Lw��=��;ob�	#e*"7�����P���]-�*����?�(��2�ÛH��B��X-]}��&dt��$� ���a9$�w����Q���-��`�����H4��~��X;�fߕ���Ͷ�"^kR���m��o'U�%��W�Y�RЛ9�}�:�3ts���mbI��J��N��,���⇉]*>�q_��x�G�3�����̻=�<�f�gÉ�G3����_ �'�E|�ך̜oL�� Xĭ�zE3[.���E0��F��S�ʉ_�	PCX�*�D�\������y�6����)�c�2xKK�ZW�����?��D�����g�g"��G�o�,6��d����.(���:�Dv���z����Q�1n�N��|�¥�p ƌ��]�ݫ��h-�z���wɳm��>[W�w����,��#~=��p�L�sO���9��&Ou-�v�"�_m����MO�+Bz:-�P� 3}Y�t���Fy֝3Ӂd��
s<&���䐲��p�%���=�W��m�1c��LQ�R3�I ��F�\��G�@þS_#Q��Tx ��_DY��`�ϣ�ܯ3�\K����rp��w��ڡ�A��f�B��"��C��NI�����'U�ETӘ�Bȱe-?��Xe\�h����_	�Ӂ��\B�7���a'���T�JFT_�^\��T�/�LK�yJ��k+d����׿�b��w�/�y��Hۦ�-�zh;��%���˽I�0a�β�Zbn����h���O0v��PO�Ǵ�(d���,� �#�,�=&�օgZnUZ7�&#O%0��vHd%|��y�"mC|h<���������l��L��y�-���\���aIr~���$ �6��<���}�f��=���g�Ge&�?&:��:�2Gd�$ �O����.�]��3��U���#ZǢ��K��/N��u�������Yȭز�7���Xb{B��^ƣL9��Y����S��$Pi���ا��� P������{-*����Y�>��6���A�P�x��b�5�u��Z�%A-Kۉ�hSb���&7d�s�.Cz��&E�3s��c{FU�Љ��ӜR����ʅ�嘮^��)��=�C�7���M�p��!��@�B�3�e�S$��������j�z~�뒋&���w�Og��rLty���@�/������0�|��]�d�F_"�@ Քή.~~�##j�w�c��U����W;.����g��t�#I�����H����]a���m���5ɷ�j]�%���r���Xي�aݱ릚*K�y��4=�gT�QZ�z����CQ}@���FA��5��7L
x�M��,Ӌ�}��
��y9�oM�͊[W1�M��Xt J��z�Mb�D�Нb��w�|��+�����[ZM</&��9��K[�ﬕi�k�3�@�<ϟ�������t{�v�� 8ޙ&�&��'.X�E���X�..�,\�������C�RF
���.���JT�����_K��Efa�vn��]�Y&	�<�TP��*��o�2�䚲[ۧ
�4ez2����׎���c��-9ju��.Ksr�n��	��O�X~ֿ�]���5���Q\�_Z<)��C��M�5׎>�������T���\PpMҽ>�, �����n����= �{&�3ms��i���ީ�����P�1>�Y����=�Y3Wa:;7��j�
& � 9��۽��@��0�7e��|�-ߥ4!��z܄�˥G��%&��k]���6Ƈf��9�-ebK㖶D~i�.&��</��.�b�1Eag��^�<����&i=W]���)�z��SC��F*L��9V�CQ��5e��3��^^l�����CB��b2���A��q��Y���hť�3Z3���$Ҋ��EӔm��TKw��G�U[_���h�?< E����OMT�=a�{�ލ4e���Φ�����*��79~'�ɾ�u�uw�"gZ~��g�kVS��y~����J�	�i½�9g�l%�-�]6_��#���24��-&*M�*�~��vrۮ{!�kv�(�V'�t
j�&f	���T�����Jƺ(��20��1_";e#��<��ӶL�̎�$����pՑ�R5���	�˂D���,v�4��Y+eoD�%�?]}�����{�z�<�%n�@��6��_YY��O��6��9�]��He�������f����������~[��_�J�	F�e��ʂ�����u@�{�3�J�T�M<��c����
������.���ELQŎ�W'��F��E�➃���E�ye����ޓ#����ː4k���?��!�>�Cv��.xk�����(k�O�=�7'E��
��8:��mV���0���,��ty.�TX�������ڰ��.Ὧ�z�V3������1�axU%	&�ጴ;:�I��+�q���dv���,���x⃪z��;�xFT���8 JT������ǞQs*�/��q���bh��;��r��k7-hЄ*�}w*
Q�Y�i���\�<�.���{�nk	�G�D�a��y��7��g!Ce��'�׍�2������J`�;,�}�P��.Z�=�����gz�#$P��o�;��^�;z?Ú"�ȉ�����8��j����㘥��,ˋ��{�O��𬋛�n�|����I�w��1K1�����,�{��4�ǧ/)Ws��7��[%����H6��{~�H����6��y�~�$�-%�l+녧�*�j�y�����uܻA6&��<Έn ��Nr~Ì��f��};����-�P��s2�04�0N�V���#e�6��G�ͺ��T�R��@��%5������4� �����$����!ͫ�����	���^7�-֖�������x� Dns�,�Q���[�HF��
_>/X���wR[�,e����t�S�ە)[!���j���<����,v*�8x�?�S^����m��]dRz<�0��-M�xV���}9,7q�~���� �X�!"��y�i��!�[^��'R�KT�N�	��r��%Z��TIyM��7~����e�ۛ���>n��+��5�p������2	a�����-�wN7��x�c��N�J.�|r�>)`M�ů���~i#U�Ej�Xׁ�󹂦�^����<i���E�o8`�2��S��d��O10�r�5��)��2æZo+��DŞ4T�w=��2J��Z��qh"���lJ�6����`�U2��q�Z�nT�ө����-���(O����~�ѧ�u���U�JaM�V�F��]=F��F��8��(7���3��g�K���̴;ߦ�.����L{d�'�R՜k��߹�ۿ���:��ƺ��_/ݤP�~t`�B��ǉ��tغ�9q�[h>yg�����z��L�`�ۿ���xo�~��)��tn�A����~�)a��ӕ��	wC��ߕQ�ǆj3�g��g������rԻ��/�4R���]rG[�{'��`�o�V��w魮��P��}����e���ϳ�*�\�oORW[G/��c?B4_e���]��;����rO+�Y*����DU��O���i���v8��<�\{�w�oFԚ�]����KƪQ(��p�6�@��fi��բ�gR{;�˥ Ih�������wu�������&A�bw[*E?~Ȕ��:�,�����l�ٛ��)7�oc�ﳨ����v*�8a��)�9aI%���?>�(qv?�|[Ԃfάk�aJ�[����~�cN�.�p��j��۫g�N?d.�a��B�*kYL�n6�9�(j5���_(�*MJ�� @w�i����,��Z�C��G��	��H�N�#Dab�g?J�,⯱�������n��ߎ��kԬ�Vq�����y~��U]<�8��qh�m�CQ M�3/(FG/�"�E�����C���޾j��`^���n��.��Eo#�	Zs�����~݁!q%.sG�+�; ��|S��������)��������L/SȒ�zF5{\��{(�i$5sT����ϰ ���F�K�_�t�����y󅦁�b	ϛY�{?��:{Rk�Pl�
x$�P���Pԣ^q۪2($K��d�]���H�"KBrr�Y�(������g�M�h|����&��N?m�����r��Q$���,<t ��dri��j�2H=P�\.���p�F�C��QLa3�*�q�����d��h +�3��^�y�r1l_��V{<�{X�����_�e����b7D�i���J��-�ꎌ_Zyف_�����Ny�"�u�8#J���T�����P���A��m�[��At�i6� 5����hV�>+_��d��TV�ta�3��l�
w�i<;���7В���v�@�lP�ca![������Pԭ�UY���G�9�zF�~�6��w����MCS&�̢ÖC�v��-�
�q��_���a�c���;$u2YP- OA��q^)Y�a���~��/�$F�^*�fNW�Թ��yL��`������gy[�7���b�|DJVwĥ��)����j�Q<MuJ5�l�R#�:%�6���˩ʦy��N��� ���~PL��� ���{qr%V�ty�D��N0י���233�i��7�R4����L���vb�I�Ǌ� �Xی4�=Lq��SZi}$c�'Z�9jc�I%̃g&���΁��tM1�v���RwB~-�xWw���]9��$�l��W���1>|m�r�6$z���c�q��!��m������Lԝ���	�s0�Aj;�
���o7�ĕ ԒGj*8ǵ�Y�xN|ʧ�4�P$ A�?�&Q�S��i�GT�5Zנ���r�h`�3�`�Xڱ�;hm�.��B���������j�U�_���?����SG,��vvz�Y�E7�%~�\�W���*�a��x�%
��=�e�E��˦҇6�Ň�ch����w��+�o�k@d��T�(1�!�F��ơ�����eM�}/�x���)ۧ�}ȣ�4�`�3M�U�Qȷ�̼���/0���e���|��bs�G
�Ozc��cʏ)T$䋕u͜qs�}����8[��nb��ܴ	���⾨���ۻ�l�R�=N���gq�R�o��/���'YrRD&�� �@���>y�4��(u�l�Ѕ�t`%�y��P��@�@
��x5�-\�?�:������>��հ׺G~��z;�_��QM}�]c��C�����������H�tK#%�%�)Jw#� - �HIIw��t	�P�C��9���/��}w��r��gf���~��9��xA��q*~�c�;�nVa#����j�M7^ͺf�3�>�|�)-
��}��#�[���9�)����<c�J����R1Y�rT]fr8ȈI��W��(�=��hHIK[j#��HO̤��������á�����ѹ.��_w�3�ԉ�;E��d�5��qw(�h��4z������_�	;�� 1xG��k=�H��']�G{�ښ_��a�;����֥g@��t!�'�s~Z�&�,/%�;ߘ  �y&�gN����V���3.�
����h�B�V�����{8��a ���&���7��
W��e��k��;}����nJ$����d�x]�z�T���߂�|�����t�Uhc]��#����!BLC���5�b�s��:,n7�b�
8��J��K$��U��G��Y���m��o�ϻ�srp��9��C��=,�1nC��W����aþe߹3g����~�h�������ɛl��O�}�[	x�W%y�4�J�D;hƆ�0�Ϗ ��/�v$����$�����9��贁g�4����v���`�������f1��"��#/�L}�Sax��έ�+KK�m�sk��є�"�N#N��5;�v�
s��szgL�^�(�l�В�}�dlde"P�hl��R����'Y���;m����'{׉S�|��@�3�f�]+V"��l��!�`�ި��-��6��؍�։U;�By�Uc �3Ky���<�w��������W6�M��C+g��w�M��o�����#đ8x�P9"��P�W��L�É��+���Z�����o�#����b$�!S�L�Y㤁:��=�y�dO�N�+�jmqmw�r�� ���r���V=3`)�ؤ�3S�e\�X���,k<=�+��
\HMD���^nx��ާ����gO�p��D��h,�?x	�-�O�(ӭ��Fl�<�Ck�e>�Eg_	��e�S,�E>g��D�
*��[����pEy%�JG~�
*�2L%��;ڟ� V�CgFd���l�Z�>�c�&��-�T����8�T�$;�(иs��Q���7KK�[��h�M�{�
�hl��!z/��.���2��Vtfn��IC( 3�,͛������O^��n$�c6�� *6���������U��k��r�#rک>J�]�>�����b%�yK++0O�x�C�;��S;�6 v��|�J�?H̿o�x>���mi��q<{�;1+<K�"Z������^:-�q;|1+���j�����+����\C�dGQ��Uζ��ӵ�<�ZN>�$��og��"�~ڋ&��Jc�y�g�g���
�L����ʰc�{�7'��-Խ:S�:F�C�%���V�o8.n�5$v7�uZL�3������k�����8�|��733������tW���P�%)(��o���Zʒ�λ��ٌt[m���n�=�ZW��10�&R�Y}�a�jA��Ӹ�0�1y~�N�
�۰o~ ֧1��=����@�!"c���mc����G�.����Kg)���鬮���&A�Xs�R��f�O�s@[�4����wh�_�ȴ�uձf
P�H��(J���z�f�k$(����<8<��Y98� �6�\����c���	C��C���!���i��_�"~�%py��s@�[��G��
�}����8����'�u�O�(
]&��`��h[��+�;��uO ��DD���H.��w�"5=�
P���؜���e:��K�\U0C�.'�F21&ڠ�Jw3lf�ݦ��:e�N�������D8S��;���D�(m��@����xؚ(��\���#s@�͍�DK7���N#^�B���H XA*�ٗ0����%�������� '3�	4������� DX���#��7�W� Z��Y[N�I}/��u<�E	3�Wk���|�Qic�Lx�B,Kt�2N�]����`K�쿹)80D6 Wz��Z����;�����h�Fɴ�Ƿꞔ��LU�E���Ȕ1`���2@�[�����s����vfV�����u�`b>deQx/1�0��P�Qh'�-��,\6��/�텓�LC�j��Y� ��	�yW=�hϗE+��1RRR����s��e�z����%RG m���Y�6"�h��%�w����jq`` ��=����.�]�����1dLҸPaξi�d�<R|#?��C� J}�'%��[S�̺5z����yMؓQ��2��kdf*����M,�[n�w��!h5Ba��,Y�n~���EӬϹ�Ҿ;]g�9g�>`D&d�|l�B����Gd�W"�;V���OSӸޥ[Ih"9�]c���@QFk����W���t����9{N"�=i�q~���/-a���t)���[��� ������V���w�������I䂹��*��'!*������;(��U�Yz[8�'�#j5�K���Oc�ܹs���-C�[������f�}%�a���D{�=qő��L����A��L6�Q�Qb:rcI�#;��Ye�sq�==��7;��ҷc����_�d�:�id�,�1z9�e�9���!������r�K��N�ʐֆ}Q���s��m�OG���!��;l/oo�������� b�rP��=ز��U:5�P_V���� ���Z��$�y��"@*��P�͝�ƀ�f#�v�׀��������˧��GT�+�r��zL׮9W��Jf�ѭ�[��y�	=9�z�EJ�J�g���jz}�E˘؋���O
D��<�*�o*����-����Kl1�w��nNHA^�i����獭#���{�d3�tI�om�
�nYmMU?h ����W찈�:�%H�E��7CԐ�]�@�X���@GC[�Q��Қ���������R����p�>���֑��h�e-��,^t:R���
�%~H�����I1O������zQ������_��{��ť��פ��[�bF�K��:k�|!{0N�yW�� ��_3Ύj��2�U�W�ˍ�ww2P=ަ ƒՍ��Yk����H�هd�k��}]p�QeIDu�R���������$!!IIJ��������ZH��>o$�n�4�ΨaMFH8��$��!��k�㓮�ׁ��9[7���Ҋ"@`��&Pz�r"�=ߨͥGRן4�����M�V_
kk5��X��<}-B�\����K0�`��tO��c��T��a^x�W���]�r0eUF��O6fye���� L:!���Jˇ
0�yW��7�C��UKݗ]�\#����z�6�]aR9��f��C-��q=��2g�Z^vEƗ��<�����~6744��n8ZT��0w�䞞��1;���v�P��ǳx����Aن��������ihm�[��C4�!pf���r��Ƹ���;%����@;[?)�������l�D�gz��e�Z$�� ����d�Jr^!@L��ƛk��˔<�,�5�	���+岦�a^�kѣ� [�1��P�Js��1��"2 �WqR��`��̟�e`��ow$�΂c i22nf�I�~=P���4�2�z�~*(wdo�������&��J��D(�\?|��A��S��jA���{

����A��.�ߓ3��lc��8��������=$TB<6�!����A먶����x���4DGGǘ�NQ="�G5�#�9ZL���@���°�#TTTB��^o\�u���R ��Ϝ5/0Ho��lN�}���v
�4�1춎>��@l�%�7���/��R4/%�ۥFVx-��qN����ùh`_@AA �cI�B�	DP5��U��+C�xg�R�$ײS�¯l
h%�*� �ڐ4�� ��6&���ނK��Gn�����<o	f����qU���=pam\/��e\�/[x-�VĜ_/���� �MO��<�].�q�p6
�Ӈ��9p>vZ��N0" 20�G� ��~�Qw��p;WL�b>H>���_�6=ƪ]�$Ϟ�#��Vh�Aܪ#�%�8<~Kt�,�t7���夤��&0��Jp��}&�x
��P�ܥ�v��f���*��0�F����yˬ׾���ӷ��j A�ٳG��=�!�\ 	�r�:�icIc+��9�~q�t�kp!�3!H O�O��7�}%���?�����6{\�ϕ�mbd�x����2�N��4�`���^�ƣ�y��<�A��A�G���2]ƙq�q*��OX�i`���Q���/e57$����
�7��GGG�j�'���MsU齏��6�ZK1}O:tZ}�?d�
l�D
��r�|��G2$/4O�
��O��#/�2���MMiT2�������0�@42�b�8���r���֮�0���|lb�Qo��ف���nG�V��5��H__;�x��Ӗ��D��O3ė����>�&��T�\�|����t�taB��7N�ԓ���nٱ26�XXX��}<<<�[�v��^�Fؚ����7�m��~9l(����"5�)hg��.�G�Z[�0ܾq���c�p��ȍ�;o�i
�yy�\j��"�~���ҽ���f5����Lz�e��Wz�O[�vD���d�8��~�ꒃ��q

꯱A�d��8��3` #��TٓGݏ���*�B?�d���2w�ϥ��nb����bn���[Pyp����~`��@�ǟ�Q�8�яQd���n''���������<��;����#�BDܲ���uZ?�88rV2|�#�����yy�� bC6��Ah�Q7˄�bE�����9�Lש����|�n���M5U�C�+zxx(�󰡱��r��(��[E����S�?�p��fJ���Gvw?�9�JK��:�z@��I�����;^��٫!���Jd�&-Lman�T\\jn�����êh�)y^s� ��^[���YÅX����zY[���+�yGtӫWZ��œ�R�	\������8~x�
���e�Օ��������/�+Q�Z۱tAO��F6�56�t��I^%�\�Iڃ%y���D��h*i���}�.�e����PSC���:���=dz Q6����*� tK���s>���HR���@M��N;��c`%j:�c���Xnƈ�>����#��z--�I��� �;��*b��2�'�#�R$��-����������x�]�
�1��+��>[��m>�-�߮�9p����h�-�ڭ��,�FW���d྄�&���i�P�b���(�����̻P��7$)6��>c�� ��@=�e��U���� v���,|��ݴ��5��x�šP��[���aK���
��!��^���c�>Jb��CK�
шߔ���H��î7��bM��� ]���ͤR���w��V��s�����:�������+�_/����-���� ����"��=�-d�A���P1��~���Gl�7���6�xg����/�`A���H����ɱ��ފE�H� A�=m�ݰ��Rp�&�UcS_�8���nЖ�n9��au�m�!�k .^�����_J���QVUN�1
.<vh7�o���Es�WYѥ��@y,� �a�E�'9`$)�O[ʀ��ή�[�@O��=�U����^`Ą�8T�uЕ��|uO��ؚk5�k9���V^^TL*'e#��a�5���Apǿ	�Oa��������5!^ޤ��">���t�t�pxo�A��3nV@ՠw�FF�x�%��;�u����Of���11����������2�7�GQ�d�G�C��U������+T��|�+/^����XZX@G/�N�6���	�.�z,'���:��EJ�7����$�z,��BC�A8<?���K3pH�9O�Ș��#	 �T�����Pۼ�VU`֘n��SeR<��ص좏zL�����������2���daz:�21@2Y��a�. pF���ƝsG��&�z߄��<NKC-����?k�^^M���M`J8�<��C_�M}?Z���+D:7�!�<����)ͱ�|C)�G\� Q�ߨa5^m���=M6� 2�c���rr��K	�_�{���;Y[�)ݶt�fYZ����gC	@'[9;4�4�� C�xyy�d�ͅ�Y������j��&B�r�:�%}�A�)��bG���R��/]RR����cL�jgg7�e~cֹ�J"v��J�Jچ�߼��V'H	�Ywi &G
�����'���e���y-���0(��wa�4�%���q��/4�8x��(HlO��7��#P�����s܋H��y��&���b�k�T�{%e�ӵ��M�sw�&��,��Ӕr��ąn]$ ,��ĵ}������R�ٳg�L+��п=F��-����n(@u�������d���]�ѸE�⩇��=�>���2@�Th�x�� ��:I��RF��,�X;���2�n;Pr%���.��wQ�.ll���J#j��)����y
,T��R:�?^��/�4 q s=@����%(Xbs��E"?���V��9Z�Fu�����Y�3��9�ctK/G!(���3��he�𒖖���#��׻tt^��ns���]Vb��T����KD,���ܪnn��C%��J7,��~��I�������2��ƿFio�X�V��oK�L�l&y�����C���g&��xy݇vD������i�l�A�&Z�2~,���� ����P����񳖺�^bku+���_9�VP�|$�-m����>��M�ޯ5㸍�f	��䏛�nF�}�)/@ό�E���$$$�VV�6�4��ٵuff����m��P��m=;;�r��1��,���ЧC)������Ȥ�� C�]�������Jo������&{2��Vxxx�)=,/��8%�IO����k�ptMeL}��f�gK�?Sq#���4�������§y%�hN66����ԣ�>O�꠴��ܳ�ć��s���g�`�lo�܌�pu�����s�<Z�-�V̇P��`��|����weeZ�i��q��g�^���B-S�,L��3i�_����#N\Pb�˖����	(��8��_~����*�,c�6)J���p��� �1�y�gg��3�ffߝ~��������؜:�������22XI�?y��j���ۍ���ө wX=�3�'`�GS�*��!	`���#��&�B��c���)�Ig�N�?(|��|�U&��,�} ��)���w�@߁b��@�X_[JᲒ�����?�*��h���9:��{�uq+�{r���>Q����BzE��������^���\U��@_�����n������{�M���y5j��8�+P�Q������@� �<��g�d1x$P�$���=xP0(��)�B_����VQ*���&
��榚��{]ݱ��Қ��ax��w�;G��"��^hm�ƫ��4u���y8=.�,m,�2_�������*���[Q��w�\��P�����VNBD���� �2Kn��]��_��U��>�F����6�E��p��i�e�EJX���|aikz����Ďì�{2ǃ��W��O�kk�����^�)(( ^Vur�|Q�P����� r��4��7cv��]�4E�?��&h�aL쥏�^3ζ�!�ݛ�m=\���Pu�qY����xJ �*�<V�N��E����HEق��f��$�{��\q+!_����*�*�����(�Rr��g�zJ�#��#�$$͋�:	��K�T�O-hN�9�nn�&^SEw#�ofdy	���
��ڝz�t��nL>X�O�E�i���6S�~���1�i��Nrڨ˹E&Ũ�_� ߀K�j�����a�<��_�6y�[bE-�!��K���*-9򂂗�B�{�τ@�����uK����\27�߷���:�2��PHH�6���S��־����G�������P�=K8���7)�����O�^Q[�ݟpI���k$HЬ�ڲ4��F�8Y>M�A���Q3��K�à���6����K���� ���%�� ����g-{����'��)��-X��3��)�W��߽>9��^�Oo����މM���z��q+<K0�9��7����3�^ٍp�0w�*���{F.��ι������ﾃ��� �/�d�c
h'ܐ̵�����s�S`��5��twx~����0M��c����!he^Fu��P.��G�ed�.� �o��r��Pu(eV$��g���4˵�ʵ�">W0A�cxxg��Qu�_��0sr���;��L�E&�b�?5IFD�-��]x��"rI�e�L�����겇���!�\�T7���HNo��o'�b>�APD��x�'������C
��w����O2M0���O�����b�2��Xߵ� ��F ��� ˈ^�퇍���LR&�[)h"c�p�l�:��5����K��ؗ$^���R�׬4`vh�� �z)"cpZ�{�T�\˺3l���
�(��X,B��o7p���7E,ۀd�e�Gl�X�M�Đ�A\nB��a�d���4����I{S�`C��]���(&kJ�y��-��Jk�����,DQ���Z�--��w���h��H���,Ӄ Rl�ЂG��6�³ #����Ng��axI��Z���N3�n����#	��F�8b����\�p���E:(o.*V��L��t��G�
}��zG���i )�A�W7=�r�0h�H�k`�x�噥"YO_�[ )d�۔n�(��S9"�ɁLhY�fYM���9��<jʔ�>g��/��˦>��'�U�K�d�S�\�8�ʰ~.-%�D���!���\=���[ )���
�����^��>�����v�?�tz��8j�Yv�id4��*oʃ���?����s�[���2xJ�/�P*�����θy�͌�]X���������;ؒ��6%jŘ�p׵Z��|�:�9���=h��'o���������κE�l������TU6.f����^щr=�ˋx�&I	�y	x�fR8/J��{�k�5��Jì�C�#��IVƔ���w��%�bc��
y�K�fӂ��I�[��ٓ�+ʌ�dnQ0��T���� ~n]��y͸f�]b�F��nuuI�e�8K͸>6#��]~jc*���c��92l����﹎w���I��&�ȯ�����n��,�E1��k{F�))� A���K?��,�PJ>��.��Q�����&@U;9��y`������1�gx.�[���ǺR���-]qz���ԁ��ԙ�欪�P��C�N�L�]���]
B޴qAte�T�XҺ��c�CN�t�&����Ƶ0����:������g���ɂ���8�E����T�j�*=�u;�R+9$$HΕ@0��+�HH�IB���Թ֚����@�c�/2�_}O�^�s:${���h(^Bۇ����||N���� �Y�ԯ��Ȝ�I�;��_�%w7잒�}�z8�?�'DE�+_,+j��2%��Q�s���Z�j��-�C�:&��ȱ��.��5J-�in��ʢ�)�'�w����P�X��R�	�}zd�Uզ�5>���+�Vѻ�c�x��;e�˼Lr�G%�,�Aᳬ�ni-���������j珘n����=1>D�{R%�4f�1�5��K�ϳj�v��|RE��Û�lB�tsS�y����j�����W.���/6��cN���Y�GK�E�;f�i�/#B6]����n������v��Q	�ѿ}�"��l}��6��A�P��H��ZJs��H�V_���l$^-��?��X��W��t�|w@�75�nFV��ωԛg|�j�`@Q$��%,&=$l$t�����S�(��u�`4]d�&�'d�G�o����q�?>�
��_TSx��g��:��=�mRp1����^D�U*����_�ñ�oM}����ΆQ6��2�����}� C0�+o�r�}NG��4m=}ve�^R����w�w�v��o}�����i����Y�X�MJ�Y;1P8��EJ���c�jsN�5���eNB�ߌm0|+�ۻ$������8�͓�?�N׻��\� �L�;��0�c���,��(�S��p|�ʜ���5`{DR��2��kԜsвZ�!~p͙t���N����'M���-'?��jrz\���D��6�����Q�����%>�]~nl$ZMM���ڹ�Th��1���p%	"�V=V���=
�,��e��0?����_~ԗ+lp�ʴ�O�O:%���Йoz�C������g��HG��)f?OuĦ4-�X63"�$� h�?!]���^�HM�FQ�m��׈e����/,`��D���KHJR��J�`�	@�]ZR��o����xz����������IvV�i��D�[����s��m�{ٴh��\!ݺ袹s�Cn��Um�sL�����+ � .//_!e�!@��&8�Ü3]w�C�ϣ43��H ����N�KHD���^ZZ�r�e���|��Q�oT���(ŅWI��kX,a&T,���&�W>�9�~�V�|�-�=44.nm�4??���rWBJ�9���5?h˴���֖���(�k��DDD��u�&�𖉡��T���*Nܟ���N�\1�<I����"����q-�r�N��p��5�;�ql2J�[O���UU�����~� 9P�%Y)g�\H�too���D��o����Nd\\\�<��B��;R�t͡�u����}�~I���z�KP|씠d(�aƚ���#$*̒�v��C^%�޴�V�q�]���9CwaI<���Q�W�X��eV77%@l����w����t�����#��8ݟ���L� �o�K^��|I	��m���6"s�>��.!�M����fRhh��R��(���x�Q��;�?n{�����p �Zfyl|<;/�N||��u����j��"�/z�*��}�)��ەr�Ya;�!JF����Y�1�Z�]��iM|�p[T�ٙ3&&�]zz$*>9;�#n�G�A��������������Ȋ
���Ĝ�\��].�^�웟.���Tb5^�a�B˥��F����{��|�Pי��ꇉ�
ntj��P�G�TT�`� KX�ß{xxd�Y"�>I��,��M}ਯ�oEHGG�+��72P�F��(F�.�/3���QZ�aqͲ������J�wd��ۜ�R|�V>���wycccr

�����%��)s�+M��ss�@��>�W~�Q;�E��H�.�e3������r�:�q��ylE�ō#ﰣ3>�A��D��*N�4���{ڄ:�ث�U�RR�===`>��r`ή���{<Zi̙���ܛ��EFb�
�����&=س>�����Tޟ�a��U�`&h�Xr6LI"*�y����Z�s�]���F���Opg�UL��C+�?�N��:��+|�q��$�"alL�<�u�"s?��{Cè��;���hWa��C�����>6���ڊ]��(w}�8��du�7�fV�O|Jg!g���qtt|����iF��Q�:,4TT^�t �I����^���M1] tyyY����Vl�S){���QRl�h��b|iz��Y�t��d�C|���1u�.=9[�Q��{���8,|���}�\4F�")!�|g�9I���)r\w����1����z
ۇr�V)�451-(N�Ho��e�kb%��K���DO�-Ĝ�xLz��׈���SE�����&����5F��j�u=������`"	&���9�f���rr����3��M��M�<��e��o~��>�� ���~�E�w�	s������+vVY��KN~��_���wqᵸ���:��;���q񮬬,��0R���C�|� >�y��r9; |7�Vo��$S$I�LPK�T�5�k-�� v��!���9@/��1�x.HsKK�g��M��jk����,,�2����3̼x�)����ɘ��d��N���m/�,����@�a���rww��Z��R���ۏ���g|�~�6���H�b����� �����[���8|�χq�J�|���S�s	<=����T�Y�dR�((���[ɥ�n��fgf�F򕤍�?<xv'1)��ɰ��7�����
6
*����C�J|���ũ`�k��W1-G�Qz!Yśaˡ�����Ŋ���K�̽���U�g>�������S��Z��_2���m�@�k���	cv��
��Ǡn+�����,.��?����>�mT9����2<İ=��;ra�jkr�wH�DK���ˀ�(���or<6�'^\\ɺ{U��4�Mz:)(ٞK'|i��
�?�����?;XM�id<�3����~����~k;�s�Se��λ���`t44H��$��$;;�)��H!&�\�DI++F(<ZZ!�|���&��{���M���{�bI���~�f�vv�j;�T��G���5�_�C�n]��to���$�l���_⣐��V��1�Z�Wg�����G��ض��U*o���
�����oj�Ѕ.�m�k1g�M�ؖ\hT"w�<ƪ�xr�!"J'B�,{y�8�q>\t�l�Kh������1����Hb��j�s�±u�9�bFe=��55���T�$�W&��e3S�{r�5��a+�����N	>@T�t�Stl�B�s3�h�z��X�﫩��Q�42��t�l=��t�^t��k��I��p�,����}�G_)��(b(�Ia�����+�+�iʞf5�&�� ���+ʅ�?Q�v��سS>>&k��|�~�M�Bmmm�P<�Vv���H�we��L'��~���s�W܊B�?�S�"
|�l�İ4���Ո(x�$���e�aw;m훰��������h̚��'���EH�����>ɗ/�"Ʉ#����\v
��KW��:BR�g�CC����F//��/P�1KOcb��z_�k��)�q���R03�k�9 m����ݲ�˯W.*���3� ��B�+�z4/`C^����}� Gh��Ej����ݓ�i�?,x�����)���D"���£�?B�Ȉ�H)����e)P��|�w�d���J��i�GB�����D���4:&&�Ouk�#saA�d��y]ؼ���(�5A��-W�����宮���p֯��Nb-��zz�� _�]]T@Q:��w��>r�8q�a]�r<�&�������P����`��+)���p��� �4'
o�������r�SG���
ç�|$	,�a4r	�uu�n�_@��8޷�iL3�=%�:j
{S='��N��PHQA�@���6���?i��������'�~��D����~K�fR�ؓ�%&C� K��\�h`���P�l�ԛ����b���P�or�G���	�̬�y�H��U���s�+!�gӾS7�9�J~n����%:::?�0�����܁h��t����G(O�}���hr4���N�q�N+����u9
r�N3���kp^l��^o`?���.K�Uc`s��+֩FED���k�ۀ-�=B{��|l���O�6p�PB+�	���I���=�GEy��<b��x��T��$��^� �!v�Y��iA�ѫCQN�]�n�	?�����6S��I��Y�-�������;ý}�E��Ǳ*��c5Q�Y�߸ێL�V'� =����5�"���`>���Ob�9]��\>�,*Z�ɗO��cm�]�:�kSQW�S^:��Sc�~�>`*�Çے�����G�	��9{�z��Y�BM�Dw��9t=��s�_�!"C��a?�i��D���ZB�k�i���R�}�m�����J�Ԅ��5��[���$0����~G\�e8���0�(1��R�0��쑉K��> n(f��}�=g����CC������-�r��������;,̍Đ"1���?�r�)_�r젓�����~m�׋�Ť�e�	�1H����~�òCRS��S8�uE�u� �{7�m��oT�\I�;!F�Y>�aV��ĝ��`���问�Ej���5{h�b��5��%%�0��@G��(���{}���S:��'~�͎b-,��UL��}�Y��_���n�����?̼��J�!~�!
��DV(�л��\�;|���"��(�����nZZ��i���H�YzYʐ�z�*��'NBt �?�Q���n:�}c�_��~��ƌ9��޾�Ty����Q�y��=��<�o�]�
xhP�O�oC=tϗ�~N����/.�CBC�T>����~߷�X�L$��"zNNN�Q�,N8:B���|o�X_��ج:Ռ�U�^�tP��Jďϱ݊�t��K�R�
������	�ne���x	��R�үY����2Z�lht����� �ɽ�
AHC���*�(0Y+Jo�!u2�0>�_J�a<(�͛5,�	%���.���;ctg>$A�'��UnZ^齆1iOt���Asp��K��q,�`�����T�m�{}j�)̜`L�f���-�=n��n7�.���j�֏��*�����9��
�YrA� ��֣�}��}�����]�8?����c�/��%O��#;�1��k�gt?!�`�EP�k�g$��f$9���h����'S-A�N˷�ẑ����Q���r��3K&''O.�T���ܳ�r�W�V���w?��&��k;H��67������M�Л�o�wo�t�p�NV����i�{NL�`�S�D�fa�s���k���^�,'��v���M��uT��HJ��L��ۙv	�P��𯫜����n!��Bmj$pB�O��鲛�����^��� �UwyWQU���sqq!]�o�;���A���ХCR��%0�Eu�>�^�;�6��HS�H�7���S�e|r�����s� �
JK�n�4���5��������z�����=�o;�,�*C���+��'���>�@�y�E6ѳ�b������^�o�i�{���-YW�˼9{6,��բ���4n�<�	����a�w�P^ٜH���v���w	-spq���g��Rt����x.
����bï�������H�Z��S�f��gcHoƘ�?GNM���r�>!Y�R���]{�.�������d�Q��ɀ����U+��u���oAÔ����1s[�ga�p��;��?)3���(X#�E�Xb�52��r��'T���T*6����v�#ԼΣw+^T�ߑ�o��N)��Y:��r|D�����*䴟�(}4l@����p�$����Y�Le:�$�ņ��_�<�E�$4�t�(���0���X����*ue��K����R���#���W$�V��<����tku������x�-�^H����Cl�\+W�h�ɝ@�G�uk*h���;x��=U��z��+,���-#g���\�J��{{zځ����Y�1^�u�n�+Q��/���߽斖�y�l�6VKOn-�6�}�s�J�	�7�M�����k�wK����Iv+"�������=t���-7at���d�%W�]TԎ����c�_���m̵��ב�o���օy>۽-�[z���֩i�z}\IH�`
���n����#�α5Q��`=�n;X�8�Ǳ���|/,����s���A�r�	ޠ|Z�W�j�1~�!��f�M�vC��5к@��[�1�d���O�WZX�|�����;52�_wH���CS�o�S�5 ����|a!��Hr�w�>�
���u䷕4-�v0l�\���~sNª��O\򧧧I��<����:��8knw��H-o��S��G��wO,i�m"<�>�s�/#+�y��}tz�v�s�/K��{�񲸸���� a�f��lc��ϵ�|���cy��q�F@L�J+��!�(��>����B��P�S���`�̬����%�C9����Ƴg�pϞ
S�d?��u쎇�5�6R�����*������� /qpۍ�- �Xئc�Y��A��e�JјV�+6v��\P��1j����`bv)pϼy�a�s)��Hk�Y{J��R.�k	3�n�`������f�zL�x|\'���&�\� �f�ߠ��-�)�N��A�~�kVC����'I�o.���Ѝ���79E���Lq�ǁ 7�ֱ����_86bGQ�����|o��
��u�w��B����9��JF�����8	\�oD����
Z�F�f｟Y�!���a�L{���e�7�,?HX|����}�B"o��*뢐�Hhϡ���˗`ʃ��Shc�uvvv����e&ddD�}�&p}�O�̼��"g-�h};"߯I��>����!238}B8w���$O�c[��q=�=�Q�2�tJ(��Mȁ�H���V�Һ��1�XDh	@�ORv�?�`"	*�e���+���-�G����#��
�E7X�Ơ���-}x�I:��&�����	^� �ң���]Lȭ48s�L�ߊ@H��p��= �\1��sQ�	��V)�/Q�U�i����BDW���.T�]6�EW��"��~#��4/����k�wy��wZL@�hs<''�u��n-C�20 /����}X�q��)��bf���>*`�r��9s-��_8K�]x��Y}�Y<((�d^X�ؑv���6`��]���4�sK�uZ�L���9��u0�@�EAJ`��w�_�?.�1�����*��[:�s-$R9C��)<{?��5Iw�H~9�Ld�t���u9���܎n����VR�R>Pz�һEo���s_��^wSt�|��pͤU�y����.$2.rrWy4Z��� ������ZQ?��������d��[�v�U��w~Y��ꞷ�ͽo,�f�?ź��'x�����?j���(Qq��bO�G�$��j���3M��yw�~���i-������)�(��,h9�E|�L?���P��zd O�*~��齅�K�.�F8��8t��e�PX'����d�T�)�����gi>�v�/��C��jU[���Π�)�8(�g'����))J��%L��K�
ls>�e�{��4Ү���r��;_:;Oy��W=6�slba=Ɵ��N�W<��@A D3t0T���|�/�%*��9n��C+��}<���uΣm_TX���Ə"��E/��l������C���g��B{l�WύZ�ba����� T]��C����48��Α�eϲ�"wsG1c2�t�?���J�K���Ç�3.��B+�FFFEE�no�e�o
�k�ó�邳KhK��4�'�<*G'&���HV�:,~�M	�7Q�H���	z��}}�ax��j���,���
�-��؇e6;V<�ݖu%$�]�*_�Љ�/'�ϫ8�����g=�W�g�B��X%�fd�Q� 
��������V��k�s�@�k5{p�ZVc�"a䪆��<�z�����HX���д<p|��D��U���_�[�q���=?�
�6JĲv�~�����1�m�� ��\-`�^n]{����z먪��_���8t�N��D���;�	E��� ���%�������{���d8{�91�\k�H��d�6SR�;'ȅ��P�5?���/"�t�+��eRg��]o�g:��Qi���;d((��R}�c՞gf�s��/��F��ӷvv6W�c������ζ�nj��	�]�i��h(�xS�'�	�����z<���"f���rbb�q��㢌���t�A�M)}}��"cc�S����6-��#"m*[�)��/oz,�e Qc"~�O����h�^���Dn"��+ �O<T���100|3X�������
�^���x����EYpa����Rr�l�\A��<���l��j���a,�(�"�t��ܟn�$4,��Ċ**G�0�腋�dߊ�����at�ׯ_�r�᎑{(����a��i+e���ݍwFB�V����]�w��8� ��EԋU^���n�� ���a�O^�qb8u]�����\���'�N�+v�H��mfL|�����n�;s0aO���Z�D;c�k�����d���'��q�j������r�8w�%/���r����P�J1����g߿��O��z�Ժ��'vc�w�@7�qǭu��ohh�a����	����������PI��t��%�������]ZIC?�MQ�9Q�|�}#<����>j������q���� �_n_O�iVW��:�?ߗ%���$\r���|���$%�)��/r��)�`�w��#4�ū,�~��@�)k# �����wm<�hN��y۩���so���䎌�J|h��z_�xq�|�O����H,
x�W�J�����סEC�_���jk\mr���ui�����W�}�.�Հ,dL7@����-z�@hA=������_��_^�,ں��o~0nxF����;���+Qh))�Z'i,^W\ ��R.Z��ԕ%�|"a�KD�� ����I�r��/0Ub�p`&�s�/үa�����U�ݨ�`�h�~��=$id��K��X 8c)�FW5���;�:��T+lll���ݎh��oF�p&#J�)�unl�y;����!.N�����2�q��=WQ �Y9�1��P$O��U���
�������zw���;�ߜ���<�X���� /l��#'ߥF'�j3d��+r����@�J;;;�c.D�+}��Z�Ϝ� ��'��<��,�[J�K4����S����6$څB���r�����y�9��Cw��y��*wQ���4.phZ�}��4��|�j�o�,|�9_h�0Z��fМ0Z5��-��9O�.��M��}P�*��RS��ø�5;����X�>���$�nc��+�~w�4LF��o�B�=�4˦a���!�%�٢�iNwB2�1���(�H�-Y�'�\���r���`��/19����Du�K����.r�?8�Cb(�<ɶ +	 ���p��u��X�W��ͧhK����������|���-)>~PE��i'j��ye��������u��m��|1u��;������i)�׈/�}�x��6���6��Y덏���������*�P��QI{;�L&=��0�ri3��T~42Z��^KIn��.M��/e��9=j�*�C4���ɝ�X���ӵ��f��8��}=�7���2D\��lm/-Q��F� ����߾�HH!��5'e�R���Ӻ�^ڢ��y�kg���rsss]{9� vi�|����-HJx��#t�R��(ȱR���+��KGo����~�ohV�d}�9ө����IJP��llN�[�aS������jj��;�a��:C���عM.l%.R3?���>�u�Y�h .=l���8O��e�Y(&��5�g�~��	%�U����,�o���IͶ�kE�Ԓ�� o�^��"��`0�X'!��[�П,x�*�id����2���܅p��G���ߨJ��!�p�[�hO��}.jv��Ƈ,n;��#<+��f2;1_2�����	�N�pb��(L������}Y�m�f? 1��V��1�n),�w�WH&�98�1��L
�A55�c:/������^��;> �����<v��@�ߗ5{��1�؁�|Ř$jQ�ޠ�D�G��!����3)��
��lQq*Q���G��h�;{��d:�̈�3���3��s5V��z�(��*�TTS�;jX�/�������L�Y�[px6Ľ>��Ո_�A��d�JBW'�@�_�������D����]vE�ϾO�A`�P���������	���a��d��MŴ��*P�yQ��|��)���Eڧs�P�m�K��}�M���n�B��(LL�
����~G(A�3u�F��NN��?=u<��A�!�|s"	1qx�IE��HOOo���]0������>7�ٲ���Ѯuu���*/j���k�Ȯm5Cd}�׹<٪v��tLL��ғ�gֱ�)����T���TWPZZ:�ĺ(�\�:$W�����)#����A�{���:�_�(��)[�#Z����Omzz{�s�*0��9~�� $HW(:AbN���9�3�Ъ/��ぱ�����0�x����\�H��.��b֑[�%�h��*��/��W
aHt�p����5�> �L̛�����Gǹ.QuW��<Q���պ�O$V����q��n��]�JG���ŗ���"��T��A���BF�7����ҡ�"�HOn�\�j	D)�i~�0ڰ��r���9��w��[��t��/V�fN's���Z�zO#?�U���g%���N���� ��
Q��KCӯ��Zw��������S���K�^yo��J�Ԕ��7��"#מ�t&[��!�+�����_[��Tr�r0����0�Z�Q��g����S��0h��0{R��`�����۷�r$R�E4o2��`�F--����-�(q��'K`�2��a���v�n�җ�P%wO������EO�� �zG�lv�;��d��/�x.V���-��Z���RY�p�ka�BT:���KZ��� F�<�%Rs��U�Ȼ���F["Bm�����|���Pv�;� fL�`�NBd^B���Ng�h��ѥ���	qT�¿�
�����p%d*~��W�e�X����ETT���z#�2��y�¶D=Ry:M�i������ܗj�Ҥ�/i��bTf-NO#�� [,�\?��������\�B�4G-���ѐ� ��O#�K�����̃����ZWY�9`� ����e#���A싧
��=�w�ݪ�7�;8��6�a;t�$K�%u)���lؖ�Y4����ǿ)�s�̓�E��[�sttt�qL�x� B��+'���.��S����'f��#s���g�YL�
'q{{ۯ���a(�5��H�Vm犺�q��n�|��^�����rH�b�z��l�u ����,��$e͵��~�]��m}���|���ɇ��x�	䰄ҳ��3t�nn�pm:�6v(P�
�І3�[7���Y�o|�e�����P�+N�� g��A��*�Vu(�b�A��hBZq(����}EH"o�G:tG>m���j��6�� ����I�����w�I %niJ���=f�t4��
d���$$!���d5�GA�n��"�Һ��M/FG��/�V�D7���:�4Ti�VP��^GwW6����F��"��+�c<lU@^�2���%��\�?�gY�4t�qeєg���=���c#@;��沐Ϗu�B�N��Pq�ũ��]�0�3���AߵX�ߗ��[GGU_�<e�������0��`���ޫ.ّ&����ַ)CP|�罴��XF�1�2d�Ǐ���T���,�L��jg<2��)�I%|Æ"�����!$����H��F�H�[��mXf+�h�b�s:�%����x��1@�N���(<8�۾�������U��0@��A�Z�:���
�q�I=�繁�����'��U;��u�)��������<~s�000�ؼ���;�u�����Z����w�ҺX&�YwVu!P}�2kl^��ɕ��6p
�yV��e{��8R��0�v3�
���d�͏��F�ER�Py�R�to6q�8��{��L��;��Yב��ʊ�����*<��~6���5���+�Z��Ax� @��Fv���\\�
	�G.=�!jx5{�h��jLC��S����$[]�����Z~���8����;���ިYe�)���e2�fA@}�Y���3,�_�ˁ �G�V�O:��r�o�v���ػc�fP��X��D�h�6���E�ѯ�tL�E�4S���7�8�E�F*��K��q/�����3J�T��8��H0�Fbe���FvbL���o�����߾�J�����Ǆ�_x�O�t�|(?\0����\N��l�+�tc|;��Zf�,~�΅���zn�cs����8$����/��v�h�X����H��"���9��f| ��8K��.�u�*�K�g�PV������Fb`�}!�a�fKvtry��F	���l���144��di{$�TK}�2�'��=����B��0���6,p�g>��KGk�f`�R'u�X-��x�>}�*H)��~��!�w7i�����O?����=k*�0�� ��d87���h<�܆F@�6+�up�R�v��0�‎:�	�m��o'��f8�qF	��l_y4>�꽂�t���o�F�Uqa�U6#3<����UGͅ�ƿ��������p�)����Փezz��o�c��~����N�OI^�!8��8ݜ������F47c'MrQ��W�{�_�`,9qg���g���V��Q:w1N������W#0�FFF��m����3��F#�G9��*
 ъհ�uXay�L�Y��s���$S����n�dz��O�aSl��	�}�m7f/���' �,�����w�TY����Ĵ�p��k���	�i��LR��n:}i��s�o�D�d�*�{R�c��O֖蚶��M��Q�͎��D���� $�g)G�~�������{�B��o�~��W��Zl3#q$�Ja24�0�Aa�!R�c�<"���S �*�P-��C��Y��b�V�J%����%�Gb�I���S���/�){#jI����}(3l�+���bR301�����;WOV�NJMOg``�^���r����p����C�я�j᜖�y	���UBi����L�W���qs����3)��M�A�s�v��J��� �-��EN}�*��`e�g~�ޣ�Tz^�i&߃k
�;N��޸���O�<cbwOz��i=��$��|�VU�O �*~�=��wǿS,s���{{��/��32HA��$$P2>�g4�� ^ۏ�e�p&?���O����}�nD�2��3B_e��o5�|��X����O=����jg��T'8�t��Kdx���HM���7`�0a��v��7QE;,!�q�هD��dD>T$P�ľD��L�y����m[-��T=6�됿ӛ��_ZQ$9��F�^���NF{a,J��Ą��I.�E5.~�	��&r_��s&{-�4���2|2t=ɖ8��3�Aڌ�9�����@2�5���8��;��_��<�+q?��!)�E�b����藄��=�Y�|���fJؒ.O�@$!X�/�"��vajBT[SUB�<�Ǌ�b�$��2?���Ʌ�U)��X���ܤ-np*Lʒvv���͆��,�!=��S]������.��|�GsVzR�m��3ާq�τ� h�����K[bѩZ�n��f e���!���aB"��Û�x�6R�
��C?��S�]���GW������j�A�$�4֮���jEA��#�F�JW_Q�YyR���9߬�4,D���V�v=M�>�=��|j��ebzZ�+~! �d"pn����ꁷ�Цe���FM�v�/=a�y1QmE��Yxxq漿a`����/|ն�/�) ���%�J����w����:�޽`c� e�r��HV���h�0����4f�_��G���1����0j�{;0%&&�/#���d�x��E�C���S��I}C�����}�#YD�����u��*� V�������i�7�q���-]S���!j�"J�
%��w}P_��<���w|]n��S�q�lB�|y�6�9��$	��7
`Et�!;Z���s:�5;b�Z�:��Q�D�����ӟ���<͓�*a���c��g�������(�h�Li��V�5�w��W��C���$�Vp�C���΄�Z����bc�N��/cj���F%C�	x�|����Y���!n?�)�+w��޸���<���42	l�J�l�AQT��k��0��ܘ�.a ���% �x������M�w�=�#�~ư���k��ڪ|���ƽ[؍qJ���� �O1Lc�T3+�K�u�ؗ:�N]��cD�umC���Xԫ��=C�\A�MD��A�_qЖRD�В�"kv���G���>>��ĩ���%�ޅX���O}�Q� �� 	�i2�n},��:di"�#Vu��dĘ'e���(1����M՜WdGGK��/?�ج�C�19����C2�����m���e	^�n5�>�x�#�$��/��wi�E��0���󋘃��?yl[�dR�[Y%����$����k.ܼ���MC�$0A\;��S�L�t��ưi[)s��M���HWPP�����U�
����KQ@�܂q�� ��l{�}:�k�"��` �����g#�@�ȑ�[]�Sԫu�c�����Œ��>&��}R��'RW)��Y5���b�]�	��C���JV?����"n,��j7��=�\5$1��Dv�&�I^K���M2F��Wv_и]"�	���2SЎ|����Ew�֜���қ�g�$�Ӹ�m�(���s{��R�ECb�/3�x�J�$F���J�����uH�u��|����j���\d��A���Y�r����8Z���J������v-�_��Rh�NPѼͤX�\���ݜm���c)3���c��;���������.ڹ��>揄>�&]٪d���FIuEm|�tL���>j��b�Ng�5��yK޸Z�#f����{���4�(1:�%���8�_����=�5���I;m
��'�P�HڋkZ�v-\�u�!4""a���Uz���:��M��#��~v���J���.6�KKt �C�\�b�H?��Ks#j�(�I�Յ��RNFF����-�Ĝ�Z�q����2�߫ݨ��Wͤ;4�+�������V��~>h7��k�Ң��r�J*6�I���1�Sn��S1�������~+�.Bm��M����S�uJ��׶�N��;����#~�.n�<������~;=��<�x��������n��.��l��c�;���y��HO/Z��UK���/J��oY����i���%�w=���7��cT������{�2�bs��]��E�Έ����@��9]�?z{��@��r����N�OŮ=�9ۂ�>��^'�uB���u^�q������Ԏ+�� �.8�*�$��o�$V���8��ʯ�NO�:�+k�hR�lB�!��~5���=7���w^�
���Qu�×^�;����e`���^`{i��%3l�n���'&�(q�am�A��6k�V$ ��8 %wn;�V�̳�����}|���Z
@�G���u�����ป�_e��x��� ��Z���t��곯�W ^X�|L��P8 0�ǫ�̙8[>_���.��Lj����ȥ�d�@=οa61OH�R��_����r��kbIK�J��;�����/����w�d`o�l"B�[qg~X��Ki.�����0@��o^8<ɫu돗���$>-�g�!LRDjXvϴ+�@	o���FI	�i�y^����xnf>7����t���V�����4z��R:[����D���6X?�!���r�ʢ/�
�ƖB�P�������vY���vP�M���9�������:����h���Q;��|�OO<�sx�dm�	�Ɨ�F�_��t�\�*>��34C�H3�w/ց���o����#�A,�]v�[���#_Y8��-qb���=>��CG�QrJ���м����{���87�w'�+NBxh��2^���l�=E�bO2�'�B�)S��un�(̽e���;��;�*�yZ�}�ϥ#Ę�n��

��O�g��cc;�8��;���Z������|��u�=N�&b��{sZ���6������Iol����Q-E%%
�-f�(�	=��Rz������|���f��=rg'E%F�~/����U��k(�ۑ�����.�&��)���9��<<��W�Y� %��8́��F�<!��%�=z�����F'S�%Jp'��K/�8�KJI��$�0��d?��*���>��S��1���s:�[���A���}��/�w��DE2�*#��Z�2���ʱ��֨�^s���[������Bl�ջ2{�	���%��l�uǂ�%���n:(�tD��������C�w%�N�z��(�ꩩ�jU���`���:p���l�|�=E�~����P�U�\�)9��Y������g0�Q�LNV�q�����W]��J��?'���ݴsS������gf��� ���y��eg�s!��/8�.����꒴6m����������Ӡ<�-�.<�p�	�;����մ6%�ڶ8Rp'm<�X���u^EŨ�$a����a�G�&U�|�C�7�2�/���x�M\�U�����é�4�Rl�On�IX,;q,�zBo,[ք̵�z�?��/��u�҈��������ޠ��^ ����%�ǒ��G���$�|�'�S�l+� �Ó9h~-���sR�?@���,�l�Mx���T2L{��Rc�9�Qy��x]��WV�Uo�H���B���hhi�2*��Z�ir;�!=sGz��RJg�.�O���;�W��l�	����y��=t(>��È�3�»w�&��BB�W����/yoc\��}��r����G��b�������N���S�P�>Z��˧�46N�?i�IR�}�R�`��Fr�6�to",�8\����?��纐=3�k���y}��*$䵗����#�Ǔ'�5�d����8���W��)ݥ���ѼSJ��aGx��Ir,ED;�����I���C��7�X�����W��.Bˮ����b����T/d��rp���t�;U|\_/���� ;A��cc`��GeR.A�ov��d�y�)vH�Fiz׽DK�D����L���i�pi:�q�ϟ?�J���yOV������2�E��T(CP�7�Z���Ozj�������Q�
 ������=M��Sݝ2Yy��]���j,�Ǐ��>�>�w�{��L�^N�nk�F.9B��= ؘ���↘�|ܶ�k��F��u'�k�V�[��f�'�$m\(��`�m<�%t���B�{03�_U&�8.��h�A�� Y�ˀv81�z�<�(���}cƺ�QZ����֤���T�yӳ��J�Td���gxcdw"VXNN��ǟ��b/�?��R{��O�ёǽQ�‍���Q� 	T�T���;(r�c���� ?Y0[.T��%��1�t��e��Hz:��QC�_��ͳ���0�wZZk�I:5���o�T�XYX`�����U���߫�t��%�GMe�Wl9^�|�5���!�����Ru7m2�)�&ks���+�Q�<t�����6�(7d�A��1�����+t�ur��m
��W;�����|�{���� ����_f�wn�}�!��/(@ڨd
�k$��()aifw{X���V� �av��xh�%m���P<����`�B�l���<���>���kk��z[�M�x��{n/8N��\\j�[�p����rb`����R7o���'|]�.X�m�nШ.]�TdMN��Vo���u�O�g>��/����4e/����q�e�_�n�|�o��R����'�Z�K�͚�򌠂�	�p4�����_��,�K ��$H���e�V��k���!����	)LԾ�U?i�hC��MU�y�
4�bׅ qppTl�L��S��.��#���Q
�_Y_+t54x�+����������5h�PHa�9�9i�󺻀��`Q6��ဖ@",���_ c7j!uss�zt��h��@"bϚ��Ӏ�N�����v�$|����O��vs2����̚�fC6C�:��\x<���s���|p�ͤ��F\LDfu2���"��P�]zHW2X�(��_I6Aw���p��ap�
�v4�|MO\'u�]H��~q6)�Ŋ!ٺ�9N}�B���O���"_)�A�n�B�.�肵}715�ݽ�h&��F��,�<���� ��9Jlr��|h�I �;n��Ov��?5�d��'� ~�DAE��M�$� '������E����� q���"H�T��c����͗o^�*��Pq��[�Io7���Up6'%���')l8'�fWSCEC6񾰰��P\�4������x���yCw𥚎}(�3��1�.�����m��I��cq�	�g��D�H�o�om�3��e��#�T���M��*��B�N4��ݯb%.��[�^WU�AH� 6C���`gi��	�s�ϝm�U�c[�A�6! L;����1��+~tC�:�J�����*Pd�? �Ԅ�>ָ���1{˯��0� +�O������B+�Tw�����\YN�髁�g����C������,������:aH��!/,.j��y���b�����I/zȌ�'�۱7M�b����%5Eǹ�ǹy��Ff�[$��>'��DҒM�o��(>��o�/��Z+I�\>K�/�O)��+ȱ�$��W{ �e�\nm8ɿ���E���T(���w��,^ ����h�I�Hgam-!Q��3���e���-,?�~g�{ f`� �Ė���o�?��Z��P��~�Ȑ��aS���bHB#F�N�^�Ȱ�L�E�.����M3LA���`��L {t�"�[B��{�(�n� 
��a�"����]H/�p5\��'�mE�L�uS0��h��`�u�BT��Ŵiٲ�r���Th�1�d�c#�pk:#�&H � E\��\�(�N>0f��?� .o�كOlVÝ;}�5"_m�q���B�ؙ�~��T�a����K�z1S�������Y���y��-�l�֋>���?8��gB�n�D+�cɀ��6iИB<J���[�w*�&dX(���z�g��U��'-��>�f2�.���"������.|����0�0k`�N�	h���ð�������MOO��٢aF�6
���ű��6E��1z|�����?M�络ɀ��O[\f�`�:ۆh9�x�Q�`�g��2�!��}N�4�F:
�:��z_ZzW�콼�yh�ye������n�Y��} +x���T �.ŶhhkG�Đt�^� ���t0->�\{�D�x%��6�@-T>���ewP�����'c�?��//I2���pt*�:���3�K2��(�{pၐY��QI$�X�{��^Ө�}^�t����211�+Ӯ�7�ɝJ>x�����J�G~����C���{A$N�жz^���`gT�cW�����χ�'��(_� �*2r���,��� d�M~��_�<W�Zuf�!kG��zR��uz��5�x�&�O�p����u��ʊ�>)2T���+~��7�� �;�1�z�2Y,(��3��4-Ez�2;!��Ͼކ`�|�Y���C�v���og9��y�s�,uaf ��;�͘c�q�\�Ď��ǂ�$��H�M�Ae�Zq�s��z�꾧���p�U��SV:$@U�쪾��[��Z��ӧ�OC��L_7r������d�����|-��?��{ÿ[�KC||p9����Z#�o�\��	w��:�XV�<�O �f:�j���&�<��L�,�
n����6��K�
+�-Bm�8lϜy���nֈ�.I@NC��;F��W_�a�E_�����dN�Wqr�8��Zq��wvb���֓L�A�mVz��C�H�������#~P�ٽS��;�cY�%��v����T*��$�מ���t��O�Io9�0��{[L�����)Pʐ�q}��������T.���M�i�k������	,����48
�$7��F��&}?��g�`�$Ӈ�N(�3���F?{#	m�&�G�Q�/��w�o�~���
��Q��Er;���1�M�$iiY*K`cm-el�d�Z`�dfG&���uG�2d�,���&�P�ĸ�_��N�Y��A\��`�̘�l����x�z5z.WDDĴI����Q�h(!iPjm�_����@l,HQx��6ĩ�g) ��W@I+)nr��Nj=?=&O�����嗕͘��H��13��0N�B��Us�K0pE�����oya *� ��#�E��N�g������M��e��{&0�H 2���i�N���S�U�fl��^��;aA����ѽZ�DzY�H&��[��h�Íd
�'� .
�R���ihh�P���p|ײ��vj���=Tl �����^�_�͖
�l��wA�>PQg�2l)�rɟv�u8���O+�އ5s�h�:�D\�2,�VE�ۭ���0�V�PN�ل����X��8�&g���iK������uu%7C����XE;Jr��?{�f}յr]=&�z�
�� /0�����W}�L6��� ��q�6~	�А�[|�P�����Jtm���Y��Z|����`�:��.WU�y����V���0�Z%��Ԩ#�\�C#7�������� �v�rc�`�{>56�ӽ��O҆5_�������塚~�|)�����vL?�^��(ϟ��>�Z�I��ٳ�IU|��I,9��%B ֊ҍ�j�ćJ���o�oNM��p"4޾5ӣ9Y�Vaē��gχ9���b��OL��k[�]�uL���n-!L��'S���HK��5�=��=�# q:yT�h4rA������r'��΍��U��l���"�8���!�����9��qN�8�kh?�+���g��K�nԔ,�O���HO_m�~D�����͛-�N��_PP�?^����d3v��y{(���}q̒���ɠ�����c&��z�4$<4�����|L�󔶷��1����2c�[��E����������t��?�қ�n޴,6�G�V-�	�P�0��q�;kI�;����~�f�`���$�Q��\��߹d^��k��K�Q�pU�kkk�\:� ��A��&	1��x�`���&���O����W�Ũq�mMf�֟b�1�(��k��z0�B|���#p�6.�_�=:�i񺠔��G�������A�6⹸����X��6>K��Z�U�K��0�֊�Qgz�&6J�lU���S�L�v\,����dIX�}��=�`������t.�YǙ�� �m
��v�F^[��<�X��Ko�]8�P�Ї�1�1T2M��o|O��1�o�=�BP'j]+��y�`7�T(��T��7qtTT`���rB��^�e�[����P:Z��ckN�_$���.7v�?�^�K��� # �*�:�㕝*����n��N)�܊���֙��I@�6/��^D�:�u��4j%g``�lz�m���!|. ���;���2PV�^�^�C
���!���>�LZOa�A�;p {����ūsJ��� �#>\�Z���PEN���u�<��×�^=�5�g�	*_�M{��^�P��C �0�?�>�Gkyɹ�fM/.Ƭ���'B����2���8����c��3�wGxd��4c>���N)��߼��� ".&����,̩��F��J��<L�"s|��f���l��N���r�_�{{{{��:5[A6p23ix�e���eq�p��w���+�,�Ep'\������A{Δ���:tt�Q�H�� �:~%�Ҏ�!��@�Ѻ��	�?'��_b��IT�N��~J�l��y.����r�B� V�2����" >�ޗ W�t*+�W����z��xC3���R��k�ߚ��A��zl(�R�l��&?�:�!�=Ի�J�'|@ť���nە�'(o)���O�K'"^[�o+'��X�65�}-~�(��@��u��/�텽��L)�O�=��8Oy�ǉ�O���I5ޖ�osLĞ���ݔ���]	@�x!N��b������Yv���"=%��f��E��jI;O@��K#���8�e�;x�p�K��ï
���+q:Yt8�@P�Г!\C��k�R� ���K����p������UW�����ٙ���f�I�uG�11(�(l�0�zyy9C����]�ϟ?zN�@S?�����>ۊ~>	����RB-O���29�����xo���akz�������F��Pk�_ �4��3�f	�qǬG�J����h��1HI�0E�4�X�L.�f�p2�G��&%'�JQ���y���=�U�jط����x]Cø���əX[��	�Ҙ��qt+!A�y��)�Dɪ�1���s�;�_~��N|EJ|^
P����j3i������Y|pLp)�g@|��~
�-�<��>*���)96�Pu8Y8�u�l��A4�׺Uh�Ʋ�g
��D�r���Դ hǭ.UqO�N�?L�;��RC������)��j�Ԑ�Ⱦ���>
"9���d�<�h<�ܱ�p7�*B�jI&�Io@�;�%�:\��$)"a�'&~�fec�6��I��y >��[���p��������H�����?�������F+�;K�	1��M?����c�: �*��?s�s $))M�0_oG�y���ǏZlcTʪ�5�(�5�Z��!�~�#eg`>bW�>Cx���/ڧ��8+˽=��g>T@tgt�h�~+(@�uT����gn�t
	�r~~b��>�u�޽�k���g!���(��^>�Y(��8��t&�<��2�D3B��jI"��W�o�u�����m�f�"��
|<::Zv϶x���j_]�I7M1%�#���ę���DY���ޢ�Y�=R�������������}�+�V=�{%I��=��������J��ᣝ��8���	���t�_�hղh�BX�fpW�[���Gm�I�3ƒ�mr��Y�U��XW����W�� ����N)׬o}��f���X�~����H�K����B�h��0$��R�W��Ot�G[�b��g���؏t�9غ��PX#2���ٗ��\�&�k�J???W�Q�4�����I%�}z���ǒ����v!�Td&���(�F!Z����..|����֑���O���X(I�/i������+�SJ��r�]�?U�wr"a'6�WN��&�H���~��	���\{"���?�����_�:�Y���Җ.����h��a{�ژ��� �y�����옓���mo�䫫)� B��խ�T�όe�>�c�a��vd������ �q��נ!��엫���8�p9DҶ�=f]�6�['8��3D�*��^��=p�/�0�to�㋥|�b%��H���pQGe)P�~���= U�dC ���<񰱱!�[���0ѵ��1��7������-��;2֠�a�ЋɆ�� >��~�A��[���T��jHv��(�c�)�&��KA)�����k$~(�����>lm��6�[����p2Ӂ?������HM.�߿���Cp>�R?�� 7�[��P˚�#��>�]�X���	Ϸ�#��/x����.ӊz�����B�߽:WA�q�aPǮ�q�bwsy<ୂvZq0F~f���'5�����c�B�����I4��?�3'JG̺�[Q�A��a	��)伥n6}ju�V��"��$�kě8S�v�0�vkk�d��?V<���M [NB�Ԋ����͉��;6�v����ǍC����71"�So�ѻw�6^��:��3�I���-�@��K��H����txq�N�sՓ3�p?������r��\/o�
`@icgg7��O���V0F���@� �P4[^_?�t�77���� �4)�����Ծ�ǽ@G{���SS��'�v^��G���.t����B�[�^�@_��|��Y����`���/F�O�Cx3�欢UG�ĥe͞��̴��WaLƢapXX�X$��Q�XNت����)&��eE�é����9���M=T���΍��Iy��`��	A���k��f�i�op�&�Jo��	��F�(qܞ�l��D�8���j�C]:Y)���f8_��L�1;+�/�0vw#�d�����Q�B��ߒ�j�t�$�����tZ�n����{{�/���ǀv"""؍i���7��͑Hp�?.��PJB�j9.`�h;��0%�7* 1GJ�J��Xsb��NƉ�����_wL���1��c�|'_&BU_���,�X֤�FMk�/"/��kt�teD񊚷\��_r�\3� )_��Y�[P0\��5�����rOc�M@�2�� �+���ߖ7G����-�_b����m6�͇��,u�(�ǂV/�����UK��
xA�ݾ3�S��7/	�̬��3zB�,��7���17� ��%��h�iu����ܼ.�:�q�{mB�~/1�@
T���HZ;�E��lt*�<����ĹOJeҴ�\�
�h�!+����=E�����Y���Y��q�sų�&����}�g	ކ܎"vz���3����jfD���5�"ʺ/B����%����d�n:���NL���:
���7����+-���-*hNB�Cpm���
^ 2F~�~����Z�������M$���q�@_'K�H�(��0b�'�Ѿ��|�΢f~rf���z��K��4[�I{���ݓ�co���\�i��!�7mkT[0��@.Ƣ�3eY�N���h)���2�n�,�ǝV�w]�b���0�	�4��`�	Q�����efv6���@l�x��C�U�Eյۡ;�Q���NAZ:E@�a@@JJ:�i)�n�����S������w/?��̙a~{=ϳ����g�U4/�t��e����6X����Ѫ"_�E�KJ�Iu�t�oP�i,�K�Ͳ��#�بʨю��^���t35d��|%~F��[��Ǖ�e���Ҏ?�B\hx3�MdoO<�!ea��)otv�u��ʧ�#;M�l;�,�K����˦�r9%���p+E6� ��1	\9+�Ayt55���o߾���_;�����T�S�9,�4��]fB.���@��Lkn���Xy ��}$�gy"�L�4�pO�of����˹�y!���Bo1��'�����JJ|��!T����#����"�o�*U��l���$�e�G���Y���,�qRĐhB���W��9{�9�@����Ê���.YG�╈],5��;;;��bәb)���?~�E��>4���,����2�ߧ��>�ub��B� ��
cXD�%�E�9�%�3��3L~<c,�	�ktʖ�(��拯��&Ya�A�vO����BV.��H7j+��[�Aʼ��O�[�,��U��ͳXmW����sk���k<����'ξ:��3O`@�`�B֛	��M<����̵H.$�"�^�*���B����rXTʹ�V-���`2&<{�/���l)#�)C��k*�_{َ�g��P �mh�N�&t�S�>��mP��@�����D`hd�82&cd4�s�}���Wx�7�䐐ɦ���i�O<�BN�����
����}i�3]��O��w�NP�W��K[�E` �'�m�M�ˍ�0�}Q{�$(	����S��)O ��Y͸A����$6˧�t�z������@�yv:�$�k�f�&�&I�j���:/����������dz7{J�����������~�i���Eq�E�\�pQ�6�ĺ ���p}��ל���û����V-d��IBA�h��Y��wc�}��؃�V����$OV5�-�2�%m$hW��C�zTQ��1�/�Pl㮛A��G����m�o�	^��^�x]���&�;"�P����X5�8�wO�!� �;CCC��rk�k��TL��r��9���].�-:�j����Z/7��R$)�@���g��U��̳|n�g1��פ����s�,�|r"��wx���*�O-�*��:�c�=[gOΐ�xUPYISm�����>���/tG��U��y�,~�0W�G|�/��*�2D&7>L�c:��lw��iQԲ&+`�\K��]y�ryE��7鯬�YW��WEAc(!ad�(�y�)f��+��`��e�Y�E��P���w���Qըh��E?Ǥ�šwR�8�>��j�E��C����X���Ag�&9�Uߟ+jC�I��z���mQ�V�I}5b��9��v{�����m�����(�go�6n���G�ńk���6���r�Ƴ|��UO��bs�Ȝw�?�/��G)4��
�b,K���o�4q	������J;5Ʀ*�����@��nft$C$i�4|w���29>Nf������5G�a����v����˩�����S5�l>��a%Vr�7��W��dr��[l6��փ5k��J$Ux˚V����߻��H���k�mʂ:8�1x��V@�N��%9�?4C~7K>��f�GV��E�PG���A5$��U~HD�����rE�FUh̛mf!Qy!"�x��IϘ���Cj�Kxr�io�!IY�ɐ��F��D�G����7��<��|m̊3�&�Ѵ1j�b|&*2фpey9���5��K^��E���h�(d��9���р���º�T����c�<�o��$�(Vy�ǘ�++y�nM�^�k��pKR*�[>Y�����Qؙ��>Bx��3�M^�J�=�+��݌�둌�z�����E��R!q��Ҍ[H��i�y����z/� �B)Nc^ � 2@�a��1��=A�(��٬,n�}<�{�����j²d&&&նUm���$����W�3�:J��c!�V��,�6�EI6㻟��X�|�J�a��::� E������6 �:2j���QF�Z����~O�?�5�3�p�mC���]�T�ݔ��Ί���gqJ�����a�އ���_��������C����k��n���P���_�KE�Ҷ6	�G�Fq��3��U&�]h���X7�5�_�ݲ�)���[9��� I�L��d��
p^Y�����!eb�I���"_Q�����,�΁#��w� Lyk�n[Lݬ[y�7F�|�|3�[��P@qL��/������&=[��_?��l`��I2E��'ě*�e�@g��;��m��m���2�K���J����!Q �����kFYN2_n�(Od}��5V�����%�Tп*��^dUc��ȭ���?LR��;�'t�����>U����NV1s�b^�9��v���������Gd0�����j��"ҙ��#z�ȇc]u��s꧗X(1�$$Zlv^�zT��:Hf����~�n�q�Ph����?Un��E�IT��m~�SG�����R����W�n��wC�K��R�q����q֓�� ���Ӕ�k*�b����������A�����qׯ������U���V���v���-)���C�v��m��>��tG2��"F�{��Rbg��:��gL�[���r ](����[�uo������Sb��/�8��r2mlKqÀ�1YT/��^�pzydTT���Wiuӳrx��P��2���>�x�nM1w�b[^Q1z�G���U�~$!'�����9�ALY_{������[�*�fKT��q���M�o�&��n��bw��{�nڲPI�|�n1��3�[�u�.���o�_ܴ2?f�d~*���[t� �D��>M/1@���B	���A>��`���*���}�A!�1��x�|5dgs�Dp@�,��������,��;�}a*'{gg3F(n���9Q�z�B�Q;|��艐�Z�e��-Y��*�T�A+P����m��Q������5����߿⦶ō.c�qc� Ѫ����}#�<*�>[���0lu�4�����٪_��./�����)Oi�ٯ���6[ﱗ�i���hDm�	m*��K�%�,�d��3�,�=��o��m�}�L�D �T�;�*�1�oa��U�����^�hZ)�� ��9�@�����-s��o��2_#q��y�1�����$�4y����{�b��0��Z�7n�x��4���<kr�v���xG�b7���"�B�/�L@>+���#���GN<�D�*Z�)�W�h��?j�8�c�233)�N��F�$�	xZ�AM3}PaH����>�b�����&I��s^);�����.輄�=�U0��y�,�ɪ� o�立��a)�Ksˌג#+uDŗC����� 6�?DZ�m�29%%��^�}�7��^�^e���t�۪YNQʒzz,����U�d�vYC.��RA6����b���  l]�	`��APdh��]�K k'����������i�y����@�sTw��%s���Y�*Ǯ�����I���f����]'@��j���߱u�M���*<��X� �!á�J���Z��HL��Ynt�(�#v
������H�f�LNM]��;�^\��{J�X����w
���}���{���cғ>wt ��Ϗ���=-����1,Z������������7�j_Mܐ?��/<��SZ��,����I��=
����7Ui�@�X��`�U9'_ �{�=yYyH�CU�8$A��76��N��4�9A}�Q�"�q���s 9̙�;�%�OwP��xz���o��]�N���Wa���A<�q����-")s�����v��g��KxO�@�V��f�B�.���Q�s#��:9���.����\�S�Aƨr����g%�������4ȵ%"����7���"3�?j����-�M���wY���y�?�IA�ʕ���苾ڇ��wkg��{+�{��I���~xs�^���~�)�e�;U;;8��:;:�V[�>z��t�<�����+������,�Xm�)GTא�����ӌ׋�qQ|��`fy!�<KA�{���@ӱ�4��"`�7\T�.$�z�T��o��|��SQ1�2�f�N����iR�_�ψ�-��͋>���H�����~0vU�QHD����-,�h� �&�<�+r�V��c.���Px�O)?}�i��*d �qk��-�p�a�V	("s�{J��'�x���kB<�:��@�5t���5��f�����<�?M��\�D!�v|��� ��a�sވ�\�/�ݑ���S4"q�P	)�j�S�N4r��0�����>bu1����~	���GA?� �sD�W}��<~���TA��z��x~�aE������� ��W���mm�$*���/��S��ކ��
 �錏��`4<�&pf�[[;�����ގ9'~�z����pm0n���W�LQ������"�61�W)/k��Բ��:��9`1,��t�D{�U*MRP�C!�k2ﲛ+��N̩q~rV���q��%�(Ѵ�d��=wtw�jrA�c�Ru��) *u�pwFS_�9avt�>��dn�?k%�������]���y�XM_m��Տ&����ϳ�WL�e:3�Y��S�ٖ���A�,t���[D��s���Kq�"���Sn�5rG��9w�ƒ��-%����K(9.Q#�O�.��D罭W��6ӕ؃L���hUV��o�n�X��$3B[�]*��=�Bܪ+mYZ�_�6�b<c�ŁRAQѪ���9��M�"����@w�v�Y&p24Z��M����!���;�bG�Ż
N��W��o��e�b�������3�MM��
3O�G�%i�K������.����z}f�r�U��0Ta_ ��U��ؓf-�Gl�c�'����l\��68���?���%v3V�l(%a�ڂyc{\NE�Ԓ��^�lp�	�Yw��f�Y���ً�l�e ����Wr60�F�i��I��M������Io�K��v`������M�`v���̇���>����_��f$;�p�T�P�1�\���jlg0q�6k��X���&�9���$X��G���Q�KEl~+0�]6�)b���j 7����hKJK���?j��z��RY�*��az�8cpgzH��޶�����Ȅ�آ���Q��*̎���I����AL	{���+>�z�}���r|���ޯ�	#7a����WĿi� ��DuD�!`�j}�B�RQ�?.U�d�@����LlΓi>��⚡�Ƃ�������y7��'�*�F� ���o��%q��? Y�o�����&5N�^]YY�z���+�:$#���,�ϸ��h����د�zߩ�M�2
�v?��+��i˼���F=	
�_}2�g�y�d�������i{�g���\���D�����;�Vػ��k�%e���on4��\)���m����Z������h��6��P)k=M� ��������Dc~QQl��"tK�̯�x���rE��>NW&oФ��2�A�Z&s"�VG�w0� ��� 8pR�AwP՞(&�ӿ��_ۤ@ÁmY��N��2::����s����5L���\u����2��QS?9��˽·S���v{?��[nv��Xgy��A��=��`d,��}$5t���jc���tt3�c���Te(p��)O+He�X�B̗�]���d0�o���a���B`1p���[&��
��V���a��R��k/UU�Z��ᤌ;�X{��e8{�1��{���DE~4�VMM�$������TyM9j�=n��ݥ�ߢX�}��\��_R�sh�ْ= 3�
���9f	��;(��Zm+q�a�m7r��ˮEp�X^\�7y�Do��5��Kuˇ���^B66�Q'��xo�}�#�͟^Cj�!��=����J?�E�o���]ۀ�#���F�I�&a��\$ع�i%��WC3������RI�5]H�e�`Q����z����kb�K=/}}y6xw�h���WSl½�,�����I��lllA���E�(>����yZ�Q~jj�1�w���,H5��f=tuj�{�v7k��h�&TH�l��'����:<×��?���y�ȯ��;�*��Y-)!
�������ТD�a�n���(0$$)�W[�T�>���=��̹�8/M=�e��8�uK�P"N{ �74~�_E2�^��l�>��!4j��|ĲR��B��z[�&��2ss�*a�K������ � ��Ms>��qok˶�E%���U�#����w�]�%��OγWVo��Rw��$�?s;�U��!���sk�����yVE*�I�����..��?
u��0U��o����2��,�����& ���uR��&ft��ԭ�����:D�	�6"d_f!Ý���ܼ�}ie2<�QgV)=���3�)$m�����G�:���&��R��C�[o|�ī�y#�SPrbp�C�����	O�R�CܺKtJ���3�3��5�����U[�4�Gؖ��(�$.h#.Ƌ̖&v�5���s:�$L�≊�N�?{�D��͹/��qy��E�����ތH'��6Ӕ�%����8�	-T����$|�Dܺ��,�����,��" e����SeU���Ln�uә���O��imjV�Ԟ8���v&{�s��x����%��;�J����L�3�����P�x�~��/C���B�&�};����C�N��US�#~���@���S����ߪ�n>�suR�gV��W��a�9E����i�i� �ҪO_噿Y�x]
�7��g �x�u]a���}�z���egwMZZ׎�"��ԏjT��s�s\�>�++t�FFV��c2��;�Z�^:����8c*�,p��S�6h��PZф�V8+q��u�j��D�i���R1��� ;v�%�c�j�����Ԧ�ȯ�T�+��.��!��[�e��ᮽ�W���An^�:����<�-fv��\�	ڗ?1�{zx8 �<�tF�w�U*V�W���h������w��X�"$��s��vٝ+n���g��jy�ʕD��FY�ZQ՞�!kt���w(6azhh�e%��
NZ�=��|AQcͣs������hF0wɐ�#	�A
�q�"�W��@Lp��*%�J��0))il֗�:��T�GjOOS��YI���y��#t��H��I�49��Oߡ{���5X�8C)��f���GR�L�w0q�E�����h���\4q�������`jj$-�/r�rT&S���u��5��A���a��x��4q�ɠ���hn��G��;�|	���7����aJ�s�����'�ݷ�@�6E�S1s�Xbm��/Y����7::��$��������,j0֜�yxP^^��n"�v@�(��wݣ$1$F�V�u�_痮6Sl��_b-n�����!/^J����0Qd�PY��_��]|�]���b
�W5�A��'I�wy��R��J�s��O7U�pcJ��q>�ӿn�B�f�I6���Q�5���\K���%�Q��Q�]��|��F�F�� ��yQ5�Mc �o��gb�����'��qk�ed�sENUY pxZ�a$���G>Q`��}ծZ�"�Ч� Xߥ��P5���q�'�p\@�k���)N���w��Q:=tx��ʶ�w�W._�Xyx��
�C�^�A�HUg?�s�$��"�Ξi�nb��KQ�]�d��"r�-��]�(9!��?'���4%q~oNĚ? ��j+��^\6Ɓ $�"S�5,b�o�r	d��i�x�H&�0��t���0�b��2Gȅ�C��%�7H��`F��6��|���}�ԟHN���ST����L9G`��G�p3X)����j�h�f��n_-((�-���0�?}�e�"�����_��x���W��ͦ蝍��n���lBi�{��qZ�݊gk���i���%��������.���33~z��6y�b�EH����=i(���c~	���t� ��i�%	�Bf��b�[�|�:���݇��t��&7���XT��[��\���(��B�ce]���J+ ƪ�N����S��2�^4�q/�޳���ظ�z���Y�a;Z��'oY�f���퉉��_���~��N��Dǖ�+��g�Ǚ���P��<R{�&v,����C�%KR�l��K�Y�a��tВei�T�����[�����wR&����!J�l+����
X��Q�*�����s�S�c����#`yy�Oi`L���R�
M����V�h�H��Ev�̢�X��!�����m��s��VkuF��	�=c|�-bu4�>�*4y�&QM��DH�>+R[����^KL"^@�Ҏ�_&���U:��G=���]�
�h"����}�O��,��q���~O��Y?4#�9�2L�f?�E���S}�T�	�é~���-���p�1�]����7�"OY�2�᮳ �dZ-
��U�� )4r�ve��!�Ѱ�?	&*/t���8�e�Z<���<�A굱�fNժ�����c��,�|���N�Y>*�-�G&Ӫ�U�y�E��W$g��0& nq�E<��e�ϐط׃�D^�K�T��k=������Y���@�r�A*�^��� �����EJ��;�Å�͊���e��}�_:!�w%�]�gr��.�l
����~T 
�����ی�H��V������'D�ǒ8�V2��!�Y��F0��bm�9��1d���Ox��3-���t�x�U�W](��>H{��*��,}�"C*S�;���.�{y�aܜ����k/H*�|���r��@�KW�9IZ�HV>�"Ǿ������TA���c�#{ۚ�A)�Y��߾Yg�B���uwU;d��M�c��[�h�*�t;�;�M�`�p���S� Y_�!pJ�@��������=*�z���;�� ����q?��nH6U�Gxnn�2�ά���
K�.,��[�T�h�z\�P̻�7��E��k
����s�H��ي1���Z�&%6~��G����x;���[��r�fw��c�ج!!tu91f��JO9��H_?�Z�-Y��|/��[��F,��1]��F.��	���P���!@���I�����n�����ÿ�b����>_���8Yɱ���u�e�]t�l�����f��9Ӳ�"�����P���p�cr����|��Qq�5r�l��{�ƞ���!��+�`�b��6���a	<ß���mf0��r�<�����Ra�t�H�8N����aF(s� }J%�Ye�����60(ׁf������cУJ\��PH��̋$��T妚����k�A�t|.��Q�h���ꕀ��pl��FO���U�f���3�4�����	0�Ҥ �>�B��$9MOG��ϟ��ҧL	Or�9��le���Y�#����3I>9�՚8�	;�����R��3G�u��Z����s��m��aɑ�	F���T���Z o�W���n��}V� ߹o#�J\�j"mk��6�%G���bG�w��J�EFXb��͛v�[@�cng߰ͲE�k	��[v�>��g�}'>�����n�O;vv�|5Q���a�$��Ɠ���RQc4�j�蒱8V��ҀQ�bj�$����4F��5ɹ���Ꞻ�)���/??#���ӧ8N�m1������~.m+��{'�O��8�a�u���M1�N����BSR�=�}�Z~G��-�nӒǓՌ3�;���tP����:��8i��#��uu�,�5�f�3r�Y �Eb7;������B�!�}��N谏Mx6�p�(-$���z�If�G��|�44D�I�@�82�px��m1$�H�Ơ׊�U��3tJ���A�Q�xbW����S6U��8ΎvZ'���o2�������L썋pth(ڬ�@7rd�Px��X����y�J�{�~���3S�:��Z���F[��O59<�;�5���?g[t��o��$S[�r��3#�9��t�>>>��W��zb��J^Sβ0�f�I�$�6�i�:���o�~�Jb��A��~!mg_ ��a�^%M�QuM��F�l	��9��R�.^�V��q+�^��:1�Y����`�z3&.�Mf��Ɨ�����^^���h��R�kܗ�gR,$������P�iƊZuՂ���`��!�
�.���z� �� ���{k�s���^���iD�k�\n�#�������h����{��
�> h���!�<��U4s����2����A7���9�}>_���
x����%����eޓ�:�v/��^D�a.�VUU���O}�0����_�Z��l��U��󋋘��?V��Fv��T��{?N�Z�`�L�<��FO�46O��·�PaT��io�=>>��T$ ������h��\?/Y;�k{q��F>��1��9=��P�eӟ�\B�cY��l�T�h=�]�L�6��ԇ����/W:�8��҇|z�\`���j����yVm��mN�G��Y�ܳ��# (=gEzK��z��z����M��9zV\�>�D�
3 ���N�%���%ϦS�Ģ�'���B�ES�8�ܬz���uu:0���G��������>��I,�/���ާ�'Q��U �jaa�J?�Eݞe2�O0ߡ	�ڗY��Ɵ�,��c�(��#%�xA���+2ss���`�&�c��P�h�(^��6$������������^)>���_���oJ�P��U�a��ˡu,��VԪ�Ǫ+l��9�V��BM��--�0ahh�r�&�o�g;ɋ;�H�~b��ΐH�~*�7/�]zf���gIp
e}����@�L�|���.�)\|�#W�o1>I ��,T��]\Dұ���0����C���v��/y���vUǴ�l�j�~��L��"ɒg�7�0���ec�;�v�+�2��F+F��G�o�m4�]� ���7�����|8ݠll�hى\%&�%�f{�+E��7��Q�N�����dݷ�z�R���2�-�A�
�T�S�(�ϟ��7u�EmY$��]>_Q�t�%Q_q%+/�⮛lu���ڀ0��%�mpe8�C�����k�E�3U޴�|������m����D��A�Pi����Q�'�������ۤj�\�����<�����
"��$̄n�(�fZ�q��2�6�S��L·�.��5`���BjZ���k �jl���o'|4`$y�� NOV��7%1��!�O��~c3℞a.� �
��)�Sⴽ���M��ܷVa�����;kt̘�p����7~����)�/�k���QK��S|%nh��dEr�����ڝ�@���cI2슸���`�FW���k�ܙ�W�>�5�w�x�9�����!�h�s�=�A��~�1w���&��)2r���~��E�=	�(y����uɐ�%*�ʊ|�XI��,�ǧ��=D˯<|�tA�������;ۼPלge�Y�ֶ��P�_�d�}��G����Rµ����[V(�&{r��U5Eؓ��o�8�.f�=,ə�}f�����	�^������i�U�+���A}"_��ns�
K鷬���N9�dQ���層�����wF�����a����U��15�<�mX��l_#t�6�{ϰg�Q!T�e�N[婶K;b�'##����٩�CT0������KnV�{B޼�L�ѐ:��r �ֿ������ݰ��H%�@���8�d�fZ�
P��+Ziܗt�� ��1Y��LG��� ��whoԕs�-}b��%��TN"W�j?nH�	�]��i�SE��~�H��ϥ�����fO�!9��q��x�0�ŗ�+�������>�U������H�ܡ5����cP
��q���lw������2ӆ�B1t�򦥥�m�������S�H)B�p����/0�}�W��	K�&̆;p����& ��a�����}��x-�����
�6��3�^
B��ė���ո0���� ���F�?���@����_iQ�M9]���T＜Bݭ�V(=�˖���4|j�-t���VS��p8��w�a߃��g�M #z^L=���aq,��l+���dw���;m;T����,������;.����a��ϑt{�fA5]_,��n�a�V=�*=�C� ��k�Z	H��Fԓ�(�~��LB߳��\N���
ߪ�~�]�|~�z������W�=Πߑ��e�]�M�~���S;[�����r����$P~�@��f#�*�s:�r0p���Dţ�3�����ʄ*�^��'[�D��N�=�WX�1_�,�y��v42�b���Ț'�Jv��7��8��/���jEV��qO����xL2.444��u������i�M�������Ɏ$��iXt�_�b�H��D..�k#�"p��&�@�F���ݼ���pM��K�����@���c�O��ԧ;�I&8����d
051��P��(�^�Lg˧_�d���1��2�yR�D2B�^'O]�ŗ�/E���GA\{�]g�>~�Yq�Y���f�|�u%���K?�tO��Ǝ������M��~������]Yht����j�v�o�ib3��!I9Py���5��W3��� J�,�:�S�E�U�,�n\K1�ӭ���=���X� m�:}�Iv�W)�]���#�@�E����ox�&����F33��&''u��K�I�+��t\�e47"Ky�˓+Y���j^EB�S���5ٓ���9@lW](��<������%j����Z���q߳���u��Ũ�ҰS�3ޏA�-����;�!��5�k�q%ǟ%���O&z.M"�.}���'�
$Z �A
��1z.��{�Ά� ��*�,Z�@� ��@G�ߧ��aYD�73�͓�)�����˝�.Yww~��nZۨ'_�[�
�j�62YL��CV�%��
��FG���źo����1�--}
�e���!O����r��E��eG���}4�z��b��zgډ_�ɑ�'��T�2H��{^|||��ٓ#_F�R��]p���/�X���#�x�x@�~卮�&3!�Ͷf!)}O{b�Wm7(✇��SR2;�<P���J|Еb�Tr�/� C�QOՇb�N�w�!�<�?� �h��^�^�ġ�sMmcK����(yh�E~��X��*3����b+̉��	�k?��P����N��P��'�'I={F���0��8��!�%F��3�跀�'�w��tٓى,D[\��[�~�ߐ��O)��*�!�h�b9>��sK��V�������y��`�y���k���8������Q�<%�)Wo[N��k�z�����=�[,�В�,,���'��,�\�m>�kO��]WHP0L�������Ϟ;��R�|����&֜?��BE[�,|��PVT�z-fx������p4d��IJ-~�#BӼ�q�n��M��i@�U�]��9����ؐ�����k������sS��������h��m�cc?��j�#����@z��j_Dސ��I�Ƅ�K��	�%Be�\�7} �,4�"FY�X[ki�ag����Xx��-]ʻ[pr/z����94����Ԛ�s�/��L��&3_����T�5_wc�n K�p�N�n���`!7��m��|������mɝp�s�����ߕĔ� I[�89�$R��
1M��ם�gR	��`�a���9ŭ)�j���|��weɋ8�-v�3_���z3��X��NNj@Bۦ���*��`��k�����
��:!E��?�@��\y��v��-�	X�-�/^O�ۿS+��=w����:*4���^&�h�St*'���ziAO��2Se����B�U!'�^g�W<+�%�.�]1��<̃}Y��#/�m0�@�U
�ȭ��q�C�2�w-0#į�ڟw���H�,�k��*�nn�n��U�n�Yf V�'P���'���AA�ԩ܂4���/p
{��\۳�����m�+ZaGd����b����F�-��"����j�'L!R�/���m��g���;ԟ��mj�O^���\b)���ﯢossCx	'O@�d%�jpߊ�,�7��5)�_{�ް�}BGw���B�(�>����{����{@E������0p���]p0v��m��s�
=���e����H ���<&�g�d0�|��%��|d���e1���ON2+���o���l��g�8ȣvŚu�17�tll|Vjq���TUUA�X��#����D}Y�`�t+K�g2�s߿�t=�2��`�������)����:b�	LT�M7D-�}��@�������AR�u��KNn��4��?�%�+��/�y"�P�Bg\�v(�7C,zЙn�dD?{�]W�R��,�PU@H�N(�cE榮 Ӊǧ��`��9-һ���2Ymk^q1Ve�Y��q�D6����rA%ٌ�Q�Pש�����,��B��5��9���^���L.��G��B���d&_����C��J�xye���S�=?����9���|N(�ǘ4��J_͋���X��j��}����w �N�����d�JFFֆ�\k�������!S�I݈���C8�76��ԣYP��`�K���:���q��#V�w��k??c���)O�LZ�ﯩ���ۗ�j�����*\�����"�e�:���a��M��|a��a��t�����2�J�v�>������Q�錰�$^�'�=@L�UV �6�Q|J
٤�0U����bS����^k��ͷ&>��P�������aIN�L934�o>�®/�:3�ɀ���J��y���+�n�hI���Y�2X�����\=��RoZ�i��"=vʫ>���g�GD3��o=:��T�|ܳ_F�q��ez5��Y�@�O�G�����B=�[���X��1��q���]�,#҅"�р�ג��6�F*���ŭYߦ���	
�@$�Q��lؓ�#�ϟ�||�X�?~KG��,\`�j^�2����>��e�c���f�P(�;�E��(�}M��h��¥o�Յ�jY�Y`*��i�<�����A��A��Xv.R�j`"�9�-`JR2n-�{�^�3L����`�\c��)�<$ ���3���n��.���5
��甙�r���%�S�4�cm:a�ԈT�iX�Ȍ/�}�f�������Ĭd$.kA ��$����o���#�n��ō0_�����3j�E{v,F�o�#���ёT��_h�>>L�6���ϊ��|v�}��<�,���{���(?�M�s}<Wv���l`��0!��v��;S\XJW�7�O�&A�>����RT+<A�
�ks0��1~1ɿO&��NV�@kU����^�a�Vl*���I@@` ���Q }y����L__��jxʾ�!��ɔ�WLտr�P�F�1�f��_1��mmlm~H>�E7�@�����$N���U�R�z����_Ljx]�����n���,�]��ʌ�J����쏙�u�Aj�*}x:"ڪu�!/��f�E@ xdh����:2��d� N��!k)����(��������}ˀ�;�w�����M���iy�c]��u_��	�ps��f���w�X���[����%�v��S��ұuT����2$�@�#0]ȹ)㣄|�&b������_���=�~G��0��+!q����{o��q�sӏ$��^�R�?J������,e�Q�T&�6+���l8��`��8l7�:W�l�ً������QM��s�@�uٺ�@}�x~umF�g}�j]P؇	n8ccbV;�v��՝�y�n_��]�Jd+�_�������KC�<,n�[߷9D��X!�B�����NK�*׀Er�y�a���ק j!q�RW�m��-O� ���ei�[�QeM"��?�U\{�����8{g������F3��@	<~<+�����?��"���ׯ�q���4d>��dRZoMܖ���t�������+_�ȿ��J���i�'v��|��<��	�E��6#`�W������D��P�e?�#�Q�f{
���w6K׏�/S/=�~��~3_�*0bM�&2k���ޞ߃�V/��"����`J�ӡX�(cN2_5&C�.�`�<<N@n*���L�=�
Č�1p�h�E�h^ݼ7Z0t*	?os�Ng��G��<��4�����I�cX�����T���3Ѽ����5@�W�"�l�Գ���ɢfϖ�xq9�ӖŰ��N�l-kO'_ ż�k�[��"U�m4��N�X��u�a������| ��(��׾�8յX�aB�G?0�$/�>�涷�&+���C���dD�T���L��c�{���@H�;]R�@��^qj�=4U:�h5�_�������g�4됅v.J������� ��o��o��#a���.��(�����b���#wgj��O�wV�⤜S��e2K[�]�`�7��a�1sZe��1g�۹&���{�)f�N|�jy����"��G^}���b3����&���C�^��lDa8k��**W�|��ު�@�`�&҉83T�k�e�,B��k=ֆFF������6F�����Ͽ��T�Ԁ���A=Y��6���o��@
��C���Gñ+·pN��8ʔ��<�_0i{w��*��㞾�!u��/�>{)���1�T��u��rrU��DU�t��wr~Θ�f����x&�{g��C�O�b�
2@?�J�0N�A�X�^��s��O�]����S��.g����*��������h��B�Y�vv�O_T��;�i������B����0R�I[�o�#C3���0�ɚ�l��n^��5�G8����8콜N���?�P��,�}�������ڸq��L�3ȻW�d�x�)�h犄���#�IDC͠�k���r��jkO� �fEt��6HU��x�M�����exl��3Д��R�@�[�a��l�-Fƌ�q��6�kHZ�s�$����l2+jXntW��n�g�da�c���	]���X��5Ԝ�NE9��s�v���6�o�(�f�x� )�O2--q��ޞӲSS����ɗd9w��7#���UK:���*��7���$����/7a�:d�Q#=u���\o�𴇦<(�щ��,OO��<�=%ȯP�;����:.ʠk�niIi�AB������{�ni	A@��K$V��������y���ta���9W̜33͹�W#֞9N[&����*E��@�8�X��Z��7%j�(+������a��ʸd`n	�̓(����nB��`|>��N��u+q{�3UR4�Õ��%�9�J�x����%!�^<�:lK�?x���(����!�� f�r��:,����o�mn��f�g���D��_�A#bQD��N7���i�y��������x�:�����b%i dzr2Pq�^c�Zf�?����Y���7|�ݩ�/����
�mk�S�þ��}!Q�*of�e�?�P@��~C�E�tۡu��E6�;	�k!j���8�ߧ���Q�g[|��!(�ZA�������s�,�w6��& ������Q����iBޗ?���~<˼��Aq� EV}0�
.�[��<���y$y��Ǿ:�#0(���� ����x�L �l~,4���?�B�bp�N���8@1���-u���5C��/0z^$O�T^�nL�o����n���E(E�����!��	���S/����}l��H���ն�☒�Η�R�N�a�WK�܁���?7�}������#����d&S�)?�,^;�0��#iC��}Y��uI/�efrF���N�NK�R7Y�l����Y^w��@����CQDm� K�6=(>[[�V��y�nӒ�h+�_�8��Ugh$�;��r � ����]9���n�����'[�_��|��U�9z1�V.�$r8p1@z��{���f�E�R��+����;�����\��lV���FxQvpH���P�V(�X��B*cGk!JW:NOU�
-�����n��?���l��Zv�R�E��%:N� �G�>�[�N������O222��b�q����
�X��ܪ�R�?��Y�
�O�ex�Q���^�3Í��\��텼��oSi�ؘ3+��)#f|�\���ڇ��,3����ղ�QbT#��@������N����AV\ύ�����Qdvf`�7�33�`7w�f�~��`���"ٳ#zE�o#�Edp��n����i师.՛�,��yu���0w��/1EhH�'�MU{B�(�<#>=w��N=����^}w	Xj��)�m�!�f�7g��~�u3�U���gY"}���U !�Tmo�>�^�{�G"ܔ鹲�p���	Q�7��I8�R�G��\��NͿ����\������"��ÿjh�ѕ��rH���vԶN!,v��������A��
��9)���.$��@h3G?AO�����2̗9[)S��c;�{!���B0,D��$���w��-�<p���`��`?�`�Mr� ҴA(G�[G�f��i��Q�vE�N��&ť�ϝSߟ{�JU6�I<� ,�Q{ɢ�,��!"̍lZX�T���ݵ�j$nVD��dLT��10e�뢐ب�pī0��_��ȳ�4���fs��&�قT��dҊ��w �G���8Hf��:�A��7sK{�F �	Ʒ�WF��M\K�Qw)A�[qB&:���v�_ld�/��Ǝ'�x�� ���u����C^ڶ(-�� rW7�r;��S��G;�#�B����DDD]��J5WaL1�cT6Z���(=M祒�e���O�cwW��P��?���q����?/�����-�����V/�fcSȊl�逩����S>�����S0�V�� +���`�q#h��o���/06��خ~�l��4H":�@x�T��K�Ѐ����ג�f� ����f�0M�}	�,nٟ�PЏ��(�����X��o�p7ѧ�P����l8�a�x1�J,���v��	�=X��Ђv��L��)����p�KFFb|�F�$���a�j�;��I�9�!qC�\۸�Qs�	[]���3�u��s�Wy��3�|���2�����s�TO�U5)���,��E��<K� �Aؕ?�&���Bq���.
pP��� ���܌>>��B�M�AE�=]�����5�
�vFʘ'ˌ��oO���¢�<�WH�VOFU��D
�
��j��\�u�Ӻ����yk1vRABj�����m��:i��2�`��j���dz_�ت��ֹ����3���ߦ|��:�r��Zcqq�)�n���?!V��M���{J(}ӭ4e�5��m�Jղ+&�,�0`H���/者<7��Z�}�0)Qۋ=���+Uc�����n>�#�6�_�tD<ś3S��#z��2�p�c��·���ד ��I9g���+���a�J�Ah���D3�7_RJ�lgJރ�S7mo�EUII�_q��
���Օ3#c@�Z��]�/b+/<�4i�X̢XSo��h�k�'�*7�Dȣ2�oZ~g���:���&��1�x��j���b���h��%�g� �5��K~[�K�G?��_KI�۬��UQ�^M�fO����f6S�&�]$��C3a�Y��{榛�}2�Eo�M0��=�a�[R:� ��dT/������l���;_?�"-�jN2��������E*l�CJF&�m-���K�Q�0ѫ�3�æ��#�TUUS��e�,~�9������x��#N���봨D/켅�|웜������&6܈��
�ML�G���>�і����T�>�Fq�z؛*ӂ�΅�K�#c}���TaOT���m��K57��$���̛���t���&��y���܁9䚨��ihW�̢���b��~����!s���I�Pr�uj���<�U��g�V�#�D��w�T��=�Vu�GC =P��pbLY3��h��,S���#lT{J,�X��%�����Ma҄�-ɖ�Ӧ+�+3��|�$՟����M�B�Exi��}4*#���d`�ZUr񦣤bs����馘�� ����K^n�����-ڈ�A �S�.���I2�3(�����loۯ��g}�.���NP׿�Y�"�����84�w�o0�"/�j���$���&���-$ue��67=���0���Wg6���e��|p�5�a�p_>f&�Wh�R,UM�X�f�cM'Erp��F��am�Г��A�XiqsíF���Ja<T��p|�T��fC]�~wU?aͮO��l����z�*���%j��hF�>~����ى,q���+��Ϗ��a�gXCf3�!�/��e~9�Dr��ˊ�D���J���M.�p�V�������α��(���3�1I�3�h�1�K]CC��3�ml��뛚���������*1C�T��s�q=�r��Ih�c� ivf����~�B����gl^�]pj*���Č��ۼ?Z�T�W��1�׽|��5��W]_Wq��������Ō����X �:<��˛*a�ozL��L�_2��fL�+ھ�Vv3f �yByjj�2+�錴:FΚ��t���|�}TXs���kǤۨ��<pf�[[0i#�/�P�8����|��o�\����Km919򨃮����-]���� 0�i<	��!yV���E-�/�H �����`�M��
�1��r��C�:q�mV����2�4QO�tś�v�\o��L���]肂.
�Iw��*�	K��S�ݒ�\jR������4��c�mK��K��>����$tY\z�jl��uX/�-HW��u���z(eнѾ�${�� z4+���II�@O�yt�GCdf�f�����º'�V��.$��w1]p��k��h/!���.C7�m��J�FO��^���G2�	�	�#�x����"�M����%+#�'���r���e�=7Vu�2B�4+�y���|�F-�X�E�"��B��d6E-�y�����u��F[�8 h{��7�~�J���E�P��sr�(��"�X6����bw��= ��F.�`���	/��[9���J����[tt�-������}w��B���li����,�ͥ�E��=��5�>Y�nM�X6��C��\B�D�udL�&�D�)F2_�-+d�����-��	<`Nm�ǲ���%8��2�;vgׯ./�g��xy��-)�d��q�{E�A��}-|b5y[�����CG��pi�rh�T�$96$N�@1�ⷚt8G�w㣢e3mWo2�+�/I0ȣʲ��̳=qmmm�k��+��S����z�	!��i\Ɨ��O�4�)"��&����-&
=�8�����(�5�)�o�X�b.T:��i��(C@��ՙ���u�E�Em�4�m���a��T�:<�܊��4�b���b�JJ:q&�E�F"	b�v�+U���J7o�:�|Ӓf��뭡�̈́���B�mY�[.�ށR[��'�Ч+ ��ɠ�Aɵ�~�\ta��H'7#��l*�Ŗ��
�� ���ύ�O~��Jc��vT.]&����M������o�FO�D�e��ߛ6��=�u�[~��=(	���-ӡ^�vm*Y��\ڟ\�i5�����'S��܆aooo,~�C>@ �}�øV�I:]y�f�1'�RrہֳO�p/d5+T���s��r����c��L��k��|o�I2��A���4wr����f��7?�ё���	�O������̜�֓?��;�M\g��a���ō�WhGL�(��I�Z�9�x��[~�vE2����O	U�B�� '��ٶ�ːP�֘�Y�?7y��r�(�ڻǬZQ"/\���?�h�Uk%�ufdf���A���A�ma��j���Aј�8]��z����~wz�O�M�!�w��o�	���"**(�&��:&��%7wp���l�����440"u�������0C��*.��B���ƥ��D�<lh�I��;U���ҋ�Zo/o��A@�Z	��G/�Y�ɞ����-���]��-7�U4g��b����/�5c��:�D�Q?)۸���oB��c�K�����$����	æ����D} &�x���6��3��v��_lҁu9H���B})����]1��©au��}:C��&�&�e��$ųM�'&'��L�ց��V�b��oqA�f;���0S�t,s������韛���VC�����:@����7�|��|�u�/Q`$�X��R.t��b�w�D�T�V��+E�*[�G/̚ϣ 9����sٙ������6E��`yl�u��S��}��D�_dE2??<���<:0Ak�#�����1_:GA:^��d�������N}s�ˋ'�ty5����0cb��`��Ľ�:N2Z</�zrv��E��㱔�	����Q�v�y��ďV��Ź�c�R�pq�\t��v�eMK"Xa�|�� lެ7��d%��wT#�CrֲG1b�8�`�����-�ջ�1�5Ir3�������f�SՅ�$�7y�	dC��f�Z/���m=n)�L���;���r�>v�����f*�g>��C�R�W*7��H`+��n��b�
��b�E����\w�����i]8���+L�i(4�T,<6�T��8,vrwg��y�)��qP��y��GG�]\�ĩ��o�./��D΅O �������St�y_����7���-$1[��H�-@]e�c�ߏ�^L2?���!7:\�S�h�Cj�mx�3Ĩf���q-��R;�f͙*�:UB�}[��gm��e�4t+�WX^��	��>0˩c��fJ-F��my�l�!M�脬22u<�z��3y0���?111�U݂%����E����/b�s�6�(h�ȼ�҇�r��p-z�+?DJR���`�0��P���Pc-��zjVf;ǹ�}�ޤ����W���i��ߨ��up0�(�[�K���dJ�Ƒ�*���)�]��D��툹���͘f3hD��̆���P�p�Z�x^���Y'!
B���n-Q���4B@��^�NՅה��"_~�������F=�������8�M���Z
񯕕�	�zz}�~��<�l��q1KR�J���z�;�Z b�C��:Uc]c���)B�:�Q[�i@<�����Qsf��꘻��;w�vn4|�M��Lu�<��3�^v�go��B2C<L���`�;���c��Pj'�8�����%��S�-������D�t��6�������֏W@B���s)()}������Z��5�C��7�^d-����'�L��Qe�9E��d�P����N��ݽ��d8a��q=�강͏�:p�ϩ=n��B�x�������-I�4����x)f}0�@�U��oTC��y�r0;���x&2��.�Y����f|��g��S�χ�#�m�ޠ֗�r����iKE>ߓw�������آH��s����c�ڪ������N�a����e6����9�����G�Un-��(1"�p��snS�x;w�2�U8�6�}��޻�f����vo�f�y�Z0ڥ�Ѷe*j���f��Խ3�B_�����{<=\Ac�J�p�"v�Ј`C�Hu��$�+>���fs6�N��.��m>sپO�w�[JI�'������!1qW:�MKh����BU��ƣ���O�^,�'s��_?V"���X��6K��M��G��l�I�!1 >M�����p�pꏹ9�ǋ��9�%"Y���c�_���d�}[۷j�VaL�t��L�.cm�Z�Z��Q������]h����_%��^�����ۤ�QUU�S�� $������q�ۻ;��A@��}%�A1�iA�<rX�oqJ)�]�V*Y�L�ܷ�_ǁ�W��+v�_)1!���F�K*�?5-��"�[,*�K���FG��Q�ՠ��2����E�ϒ������܅W&����ִ���m\������ￆ��5��Z�"���Ͱt^j�_h������a����6��ʣ�O��JK��,G��Xg,08z�G���:RU?d�	n=�L�Z���!S|��ZC��!�ښ�w��
����D��֨��κ�Yڋ��ۓص�Eiq�G��X��pv��I*}ܽM�Z�rh�WFU�f(N�\r��:�c���8ߜ�>�X�g^� ��_����h)r��f��i �i�yt}��l2�ܪ�̹�B����դTѱ�u� ��J	.��� cLA�H7�M��B��嵉�IQ=a�nr��,�H$^D6�.�	��Pf��h�y������z=�:w��S;�w�~,N䱉�^_AQ1}D޷8D�þ�60,S�4��~���R^!E%� _���C�7��o�ܤ�b�Wq�����U^� Y �,�ￖ�9]��
�A�˧�@O ��D�&r��9����p��;���n������X\��8����@��燐N��=��@�zďZ�J�[�A|n�HN\���@��8���I,>O���vJ&Z�X�I��=��7/�(9��'o�gN�׍%�Q�G�_]���uT�~|�'���Ϗ\^^��bv6�勛��w����HiY��J���*��PAK aA	�cJ�����(�� �$���2$�/�`H�緵���L�X~=�	���; ����ē�c�8.+_���9�G�&[ȣ�S�h���m��׋�x)�����.��UN<o`p�LZ96	oD���̜�;��{u����v�.UI�!v9�A�����D�,7x\�Y��2� ���f3[�ǪD�{x����_�����>#����/A\�����.���O �"E/��ˍ���*�W_{�GT���f(�������:cJ<��֪e+$�,�ZD��.�Ӊ�Nz�qq����0����%;c<�O-@�~e�c���=���A�]Ψ9��M�n���{e��p�&7�����>��U����~�j����%z��].=;۬�L�*AԾ�s2S�����~��9�awʉ?G��"??'��ѷ��X�]�-���_A��o3��W�.e)		��W|kC&���m���f��xr>]|Xă��=��2ŬO���+ǰ�L�RT-�e����	��lN�e<q�SSS{���e����
s�����7�L�jtt���.�;d�7U�U���}}$	�G�+��2�K�['r3b9�o�Æ�v=?�AG��]�+_Z�wAإJ@!�>�@�|�y���?S�9���L�s/%]ќH�B�-���"��0�\�t�h�%�'xb�_�j\����~Kl���:Jء�n����b���ڻ�?����~ ���;�d@�O�5�D��Ӊ��b��H��N����?:��Q��(J���0��LU���S� 
��=ٹSd��qJճZe2
xQ O�A]���v�M�)\C��G8$<��Ǻ~V..���Ο�C�LU�nTs3��b��F	�b/�yq0��Zfg���y�m)�EQ�Pޓ�I#��H ��V����\�ƈ�����v\ ���np�����ˮ7O܄���kik�QMOO�R���]�ʲ���w9 M�a����w��������3Rѧ����a�<��@��G���R>v�$1�+���g�^�]�D���S��}��
��(�\��Q�������&i���O8 §N.ܝ�V�zl�]E�Lx?S!-:y�.��P�9���(�G3�=.1ymaȂ2QQ�̄��>���!���rڪ]��W���BΒ?HѶB/*�h�!i��"�Яy��FSW������24���%u�#IC�\������I/vp��T�p��-���}A���soh�'�ӗ���_��59������z#�[�P���1�y�)��^a�=ӯ�v�G�ѐ�:���yP���i�b��{��ə7 ޘ(U ����;��ݢ��$���m���p���OSN��Dm!M8ddc���]�#i��c�[��aW����f*���r܋\{�O���SUK#��&G��9G�	080/�R��0�vpAEy�B�3l������Pu��/���WS�+�ej��]�`Q\�X*֊�	0B侇�s��L��s-����,������ /M~w�>�^��i��ݕ��t9 M�de�]T[XXp P}S��	٠��r���G��O	cd;��&7�г� �7и�(�u�_ʌ�v��ĳ�fnm��n�H��.�<宒��L~��;��������A�'\�W冭n/�7�$ဨ�񃀑 3Y�=�*Afe�>T�+�����bx<�s��ȶ����HICt�r��� �\|�kb3|ťh��m\�����WXI��
�.A�A�K��1��j:�Ԩ^Y<!R�*�C[�S�4ih�6��@��|�܀L��}bUz���!c�W���I[\�V��M�K�j�|�h�oA�>�L�����)靁 �Sc ���#�>����2y�3�;/�;�v&�]��)^ZڅMW���I��<~{2�i��,ysU�1�+� =��v���QG`�ķTu�G6��uf�b�@�M>��Y�2�疵�3��A���J�Gq$��YS�]�j�]��J5h ^��d���\Cp��)Ň�E���.�@	��%|r�l1&�N��Ï�B-�?J�.�m4-ol$â�3R�q��{Ϥv:m�����b�,�mX����\�PA I��K�d��`�%޸�U��6�`������F�쫵��n#Z�#���|tZ�BS�S�T��Z�l�}F���׮�dac�s+��o~��z�5�j�L�A������?�,��rkl0ᾙ�OʢQt�p4���۫&"_pƘ>�atlYE��Fg���Fլ����,|���\h�S���fI��k\W�����/�7��P�N�)��`p�����0ɂ�lB�U\m��������ؘ�+�p�>_��9�)��	�K��)A��(��d��_ul0ZR�K�X����7'I1��Dk�S�zK�?.�V��9;t
}3�<Dk��*��t�J($��X��%'*���m$
�N����.@|w�b^ �omi�����s1T&����y���3�!��I^n�0k\�uX���`:??7m�䒣s�����G�J���E�0T�5�J��nRM�w��8�����������ձ\��i��U���Ao/����JIF5�-B����.��q�zÂ����%ݺ����ِ�t a�ĩL�o��o���� _�½!��2)��������᎒�(�vL)���Gi���r�[�������������������������	���6Ϸ:::�K�l�Th��Ri�Ir����bœ��1�����Qs]�Y�8%���<�߰���qPJ�(%9u^��y��\y��S1�)�'Ա�8��q�}�r��$�L ?= ���T#ן�J�<D9l)	H�i�oArf��t�\�K���
��X'����~gN����f�vT�������͝WZ*��*)O#�3ʻ�7�G��ZDD��Ieǅ�`���6~�<`K������L��N2�hs�I�?������	}�&���1F�u�t�(��B�x��0���J��r��0�,���K�K�.�������|�ikm����ؐ݌/�
��%�6�]��kE�4�Mn5"�Q��;x�(�pVT����"����p��j.�ـ�I\����E��L��F�k��o0WO^>��F�H^��#y��cj�c;:==���Y����\���l�w~�%'?���E�FEú4D�I�w��Z�/.�,9�$�+M��ҁ S<A-�Oq-�1���(
Ó��T�@�	����#/���Dc0��S�����uGlׅx�B�xm`�'��O�-zP����H���^O�A��g�j�,�Ᾱ�y�q��_t6�u?�������/ZX/)�|��]·܌��㝚o0�*x�85[MB��	C��5t}�}�^��E���C��R�����gx��۔�S$�vke��U�pÜiH�/�p��滴	gW\շ�d�t�Jqr�|����C�8�ˢ�{�+��9�Avm��ܼ����R蓉�h��]t���w�G��V������ �#YF�C�}��շ�9?t��m�p�u����)���ȱ�}��?�ތ��Ye1N�����t��r����Ȉ��ac1$�nD�C������n�dp��}@o�ˀ�3bi�l�f�:�O�'�[�Q#l�Y)��3��Z����fU�=��c�v9�M9�c��3G�)��n�� ���GIR]���C���Ӄq&��5,ދi����nh�0f��ix�F�M�lɕ__���>�rI죲�z�Df�%W��Y�퍩�@ <rMK~@>9yh>3&g��̓_�v������G� ��K�,<|;䀒]�{|�k&B ~�
Md0[��_�_O+h0�L̹�� ߅c�+���p���c��Z�}Me�⃛@�O0�3�~��4�C,�׿�䦶���c����]�~!@�3NK�X���J��)�_	y�!)��Ī1��W~���/Ȟ� ����V���j/0w�������*g�]�:��!�'�g�f
D�O��@)~������ҙ\Z�U�Y����Y8&���U7���@+*x�ٵ��
Zp��v=n�������z��\���Qe�^��j�FFF��M�� ���Us6M���ʚ�i�Ӹc|���63��s?t�|}|W�.#�sێ?���)k�..8G���X�G�c�[�{��v|���������F)"B���ji9��*�R�^�i�D��f3��KȮ��MMMʹ�%d`p�`D~@�|(s��+s�tY�!U�SK�,	�JB.M�^�1/\ɲI(V����d��:Æ��ga�pʭ���xm>@"UU9x�
��lTҧ���@ Z����066��v!{sjEW���������/������5սXRr�F)+; ���m���o+�t3��J�b ������H��0|��ȓ�R`b�0j.?{��^RQ1��L9��/�u���!��駵	ؤ�pl{&�[A�ӟd��JM��z����{��f�-�/��6&���5�=l\��>�ᑭ�k׌CLl��ğ�_:�k`@�vA- �������N(XvD6-��?�&v�+����G{Ͻ������,�w��KN���nnnK+�@���zWW�l��v�8��Xh�uh]�*�2�"qܙ�LNI1�727G�k�&u�2���jY��!���)hS���߮,�%��p%��J�:�;��������R�κ�hV�v�1�1�ې{��`��7-�Q�R�a.)���)-m���w��ܔ-��]��>[JTmd"���[&��ʊ��̻��.�bE�k�#��0�#���8�����U�X`9�7U�E������f�I:��~�Yޒ�lb�iT���T�%W��]t=q%��ף]��$e��E�rL��ih����d���}*I��[]]�,b����j__S���7��}��'y�Ғ�䗕Y����O	�G�jz/0h�Kݢ�w�n&�l;M��~���[�8�[�f��ʋ�#�ذ�?�xy%w4�t>��A�*���� a����'|ԲϚ�l�;�-�_�F�s��f�R�P-��-%�7d	�̈́�Bƙ�(i!�;I��="��m��8и6��(�h@s�`EV�"+���)��mg���p%�k��r*}���
�J���;<䆛�i�M� ��~��O"ek�{�4����qQ���
s0�(ÞF0�A---�1�\i��{MY?EC�b��ݾ�?����3痗t�ud�S+��}j���\h0��>�����_6�C�໿�1<u&$$, #�P�����ֶ_�wQ�{t���X~I��qi���, �#��;�I1��}��y*!4n�0Ѯ\����ͯ��&*���PC�goo���頦��S7ڴ,i))�O\��@���Ҳ`�.�$F����띹�����{��dzlC�_��s�&.����Mq�jCb���	�\[�"�9�R���ӵ��&���2W/ߡ5'mr(( ;��K,��y{��g�cm��6;����)L3��~���k{^��E;��J2T�#��Կ`H�$"�^��vGp��ow
V�F��1�j���_���nT)o��3 �'w��C?��].��	p:���+z�������3�#��������"�	�i��v� ݠ���s-�:�sq_�L3T:{C���_m��3TӶ��40����6�� \@d$��{~Gy&���C��{Se��4O%����#�?�`��}��f*f�!:I�Z�}���鸊�摑��<ZT��G@ �6;��2?��i�M��kl\%�X>6d�l���t�8"+ЩjX��/ �V�)�\��q�o�o&{Δ��h��N����_v��<?���׿�i�<�M6�;���;�\NX��_��PٳZ�[��hJ�M�e�¦
7�;�2vh흰#�L�K8tJJ�]M0�{���Od���u���e����dƄquqYI�ȑݿa&@ H�OL[~>�B���o��B�!��8��e����h�J���)�N��K�灶���StT4���:��aj��9!��*�6�{	Aw�32H`D_c���9��:���j\�l:5W����(�N��n��qGGG�����+�B�b{' g��3��a��#�^�B�����@��o>�ЃζF�*�x2�xE����=�#�����x} ơY��,���uV|��	嵔
���6�NA��N�?�gy�������i� ξ0���eA�v�����W�O��/xQV��A���>"�=p:��
	��y�)?�(ι鮭��C����!����3�~�X����֯���רڽD&R3�hMI��>�»�y��v�o�9�V'�ҔeD�|���4�&K���3�l>�nGwG?��ĸHa�� �O�� ��־7B�s"�1�,R�"�G�77��F�B>���4�����fx��� I���&w����`�_k�gj�۽�tFPPw���`��Ǐ��_���|}}��)�����o���>�V��3�Q����.�?U���q�R99�Ţ�M�6�%P�n�+����,--�N��![�N�?�ᶺ�t>��񅆅�` ��ͨ��{��i�{PaЦgsɡȎ����z#�&+e�L�ˤ��F����۱���ܥ���_���8��J͈��+�6�����O�����un���G;���<���0�)��U'ſ�"���n,�xA�h���P$�i����b�SC�]d���V��qP$��9l�;Ƞ�Iæ?��O��p����rr%�������^a�t��BGZ�N��^��L��f:.��e���0��L%lC�J@1�Vj��Nuai�Z^n��܎w�!���Κ�?0Z�u�@�.���.���g!R�3Qǝ�Ke:,��5^:��$��(�Q��F؆O�3����l]G��oyV�[ZH�� nN�`-��\lu/���'�f�I���Z����������N�7}���B��R)��s�t��#��v]b����N,?�����c�:�g0�%0��Gb�u�п�ͭ~��ը�L�S9C|���pv��Q}\�\Pw��]`A�wS48�giJ:M�b'�N_#�׷ۂ�1��L��U���� ���g�u�Lf���Ps�#C���n�BLlƙ��[��P��g�zs&��z�Y�[#�H���B*ŨF��Q�|�c;We�r���DO�Cy��x3H#+������AЎTT\L)�t�5Hԛʢ�0��8��<)�`���Z=:Y\RR0���jR�� ��ړ�U����Z�sK��`�x�!Z��ëI�Sv�uz��rp���J0�X�W���WVQ���� �-̆SPZ�V^^�Ns�1�l` ��O�*A
�M��b�}�ƈ�^�����ӏ�Ŀ&J�䇼
/�E�L%@Ps��4~VBP�pu�����3���Rl��u���]���r��0E?�m�JǑc%4mo�r�}3��^��e�A�[�E�+��W�#̼����J�d~�k��/��������H�X� P=r s0�yUU�ִ)������ɨ	��9wT����]GHII)�&�y=AE�!�ٚ/'�"d�P�[��n���vZ�0�0]�)^e��}�hAA�5tY^����1�wU�����ZX�pq�����|�k;�*ho�����fNV|4�T	��B'��ZS<`�u�Q�x�t�&�+�4ц�x\#��/����^��zкR�d^s3ߪ�����3G���,�Zr"$(d����xe����5���^�݊S3n���Am+&�[sM�19"�}�� �!���e�/�C���Zx�/����М��ta܇1��{������ �CCyH����;lH8-2q��u��
���[m)]b�)���Q����M ���#P2�#Q�wك68��D�ϥ���*	���_C�д���[j �y_WW�5/�x�@dR��b��� �}_y�R�OG8=tt,LL����כ����I���p$���i�a#���P^!���Ғ� ��_�2��`^�А&�-f�ｽ.��+筕�T��-MbM�L���KY[3�2w�H�A�ϕf'ҫ;�� ��M��l�wo ����o}�Z�X�G�tv
z���H��ʀ�O4�h��T�� ҌG%�r*c�ܼ��RRRo��GG�Vj\�z�ׇ`n�6�n�`�k����, h[T�xlqNk��g�����{�4���!wB��y�!�0R~�Fy�}@`(q��G���3A�lNK�����Lhh��g}�đ_�S�11��?WR5�i=??�,WD�:�uO9��;��D��a��:�̹H�O��!��H�b`��H��(�@lu�Ȳ꛷�kk�K���ͻy:�ㆇe�45-�[�9���޼��g��q��r�.����������$����w�W�<�_�*��
ev�0����b�'��� e<�[��w�ᠷu���`@����@����\baV�lmYܠ�R3�%��#ha��ֺ/�������	^�G!��	Y�l����D�;~�_�i��\�#���� ��qeM�q�Ր-�K��ph�>�T���v��p"D�����e���}1�*zm59�@X [��AS(Xm���J���*�.��tl��]�5�n;͗x��y	Ŀ<`l��#�e) G;�2!=8�D�0�8ർ����q�ߎ�p^�R:�T�����d�x���h�kE:pa���L��q��� ~z���D��'*�?��ħ'CJ;s�O����َ�ڈ�J�m5�I\~�k����Y�&�<�q����VT�,
�h���[�Ǝ�!��ss��\o[��u.����2�һ�P2��ޜ%�7!�+ �����GW�KjqM��6A��^o�|)Y`m�i
�a�L����V�M�0 i������X��{�0�K M�LsqEN��l?�9y�����n&wn[�@��
�wKa �������V��O#��\���4�leV;������<�D�����y�F�[6QYS3���q�>
V>l�C�N�����Q��Dr��i��7yqԂoë�;�����z,,,��a����l�g�^%� ����GG��z7�J�����r�/H5��QM0�Zɀ駪�:�!�;�708�D��4^�,�K�J�i>���J����+ʹ�3��3��KM.�������hZ�0��/Y���zvzG���Hچ����ԟHql'>���ڒ���^^^�a�ܳJ�����ӗR*������zuQ'�W|�3�wU&:_�%^����|�vT��.�;m ��a��_��er)g�nnnZ�ۇ-�rv����e��l"���m��^ER��(�$�(���jG���hY�Tn8��B7�w��]z����Λ��t,@����Ay��·i3k�ɟg�Э�f�~ �e�d��,Qy���.�e���n�Ly0@��]��:�Ȫ�:%.Z`��t��&щ3M/(�b���1��;)����E�d�D��e��F�V��{`~�̈��G��f��s���_�*#�q�n�m/����lbܦ�iAT��y~yG\��]R���\���5� �;�ٿ�o��� :�fhiҰWf��K�vvf�ZP�kb8��vH>�]��0��4l��-=�HNM��T�<K��p�3��i7�S��1~�w�[��`�cx�0��"��>C���-��U����QM|���4�WB��~I"gM�;��n\�S�~����
�8�����m��\��C� !H������-x���{��5����������֚E��g���ޟTUW�����-;44PSS3q0�t��:jv�Ò����r�1؆���I�oi3��Ʋ !�Z�2"8��>hll,hg�����p���G�����Z�AQ����Ϸ�T<8��}�P�1=��&(x��r�{�u�MC�>Q���)����XYm}�e��״��`� ����l=�H��m�7{��_bp��C�A��x� �tS�׍b?r��5V���-�Z_(�Z#�}�5��9�$M��h>�+�L�)yN]���l~$�YmT��T��+հ1?@p��
o�g��M�
O���|������s������QdT���~����ݐ�g�=BL�.�~}�C�Ռͫ��0Ǡ̌�͕����rK3�66J� �
��cM\�Q�,G�oH>Ȑ#���#e�D��̬ۨ���@�Ȅ�q=�5P�!�)�p���8�;�6�k�!�oM���r��$54p���S|�ڛ�����f�SH1�:D{ �[�t��Y��u���Q�e����c�����vij+�Cc�wT>�bi�VZ*5}��;�C�RI�!S���_,��𚆧��4�@��UȠ�����*�l E:ͯ�aŃ�u��ʴ`�蠸���m���ƒj�����qg͉���0"�g%�S��?E�ި�2i!��Tٮ
/9��~��S��ښ��8�Dc�_4�w�E�4�A��+ǃ�g�ப�an�;�L�$��d��r����+H/֢m�.'�$��	dn��ݽ������v�����XT �P�A�r��}�֯ϴ
bk��*���*GT� E��ߐ�~5�i?O��������r�0c�tȞ/@<�RR���0O�9}�����|��#J�ғ�+�TP+�z���)M>���T�}���#i����_s$��Z�i �d�uT7�-E &�m?�"�V����(�?<�~�|��mp�%<�^��^x'� c�C�|KY����>&
B��Lq�Kʤ����#�/�����Y�9�4Quuu�22T�G
�߾��5Z\L��@;�m���-��I�+""�$*��B z��Lq`���냺�7����&�2O?�p����L����o%I�:I��Â�"�Gl{�+3��i��CzPQQ�u�E����*Z����&���Ĝ�8����\/G�'�0{�����y͔�D��a�	���T��}������_����a��<����H37 Juk��.gזe�ۻس�+ͪ4!4v�PǸ3������.T5ӟ\会,	���v�V	�rܯlǦ�������h�G�ϳE*5_.���Z����� ��u��hB��3���?� ��k5����*��?d����L�Ĉ��Wu�S̻�>(�/=T�pM���T ��\^��j��{��Nvmj~K��~���~b[]��ݰ�#�����fN\���I�6a%���UQ��k�ֲ �j�o~�{߄����1�ɫ$J	�%vy�J���i2�tu�QT�������o�]7�uv���s�r���gl�������]�����xb�珨���:�ٝO3<~z$^a�Rmil�n�1�Ǚ�u�c�e"-m�G���	�⧻�l��U�5s}�fk�9�� ��~�8�����Si��F577�D�Y�	�߽�0�덭*��t��_�*����S��C5���bRܥ0!���Fi<:���9�����+�1��2��͢dj|��)ͤf���l�f Gd��r�>����L�F��'o~g�=[�c�I���!�zx���п��^[_'����XxHϵ����2���ľo���ZҺ����m߿O��Rݾ�c̺\U�вg�����|jHf� ���ed*�ǺjQ]���'�q*��`��RQ�#d����p���#��# ��ZZ����muF9��P4���YX�MLh�N��u�YYY��_o4�لS&E�^)p0�l����N�ò��8��S�kd��d��}{���쵁���*�u���F���Ʃ�;2�#`B?7w
N���QS	))8@#:R���|i�Q��o�|�)�O�~u�_Ad�x'��`�r�Ntr"lY��L�(7@�b�"Rh})�C���FDn,����ov��w�|p�ܲ�.:��?�"9��a!5��=�������<����U�o���m�M&�zeee*0���,�,��]ʊ�xQ�#���Br�x�_罦f�,uB������R���G���='CCCʽ��l���H;��!�4 ?W{佉;T����>�l�m����Bmm�ݖ
��Q�Jݽn����ۊ{ɮ�o=�� �O�Q��u��6$�v���o���xI~,EҺ�Cv�\^�njj
Z��<�Wڽy�����5?�U�� ��yF�膑V�;��\�Y����7^����~qt����kY�Oՙ���+H���"Z�`H�2�MHL� ��楖X��*��5a���Y�0L@�c��.�YP�x����\�D�֯��|F��|�(�U9�o�f]R�pg-�M�~ �1��!PYl�������}°kj���� ��ų+I�`L�8��C�5��f���c��t����g@(��ңM/���uI�������R��H ����M2Nv��}�ڌƧ��ϣ���ʫ�@����"}������2���ީ
i�´�a|�=�Z� 9���oafX9d��LI,����f;�K�����ǛM���*{q�9 =���xnoh�s����QS���D¢�"zF��R���H�U�iEm\���O��G?f됿;���$�xY��b~O:i�AG���|ú��{���4�x�Ȼ��q��U�0.A��Nm���}}}��=sɟsé� ena� HU�������}�i�يͱ�l��>�9-н��3�B��w��+	�eb(�{XuA\�v�92��3�0�~Jɢof�t���Y�v<����	�Z��sm1�qT����eͥ��l�(.���ێ�����n��*���T;�b�''gѹ��+�f�gƷ��.��}�frb�GYU5�ʌwO�]����z1*<..�+����o޼�������l%Ad ��Ʃ�U��c�F?��@��}�=���W��|�5=a#�����91�����V�J^r[W�����Mdi=A����'" +����f``���� ��j���x.�V���*���>G���A���{l�X��nǔ�qV�c�t�3|i�S�w<�S��-C�ܲm$G�������5׮�!9�6=�$��:��.}Quu���2LTxv!�h 3�&�L��p21IjiB�i�0K�ަ����/�jO8���R�{�� }����-�e�BS����°�$q3v�BEJ����C݌)α�;Y@:�tGRM�`��p����y�s�5(&�%(urZ�qd�/5�" ���h+�Ã8ν�=��B}�L��8��<	�m���B�wz��f��pr�в��@��[��͛���n 9]\��b���C7d?�83/���E���׸�[.�l���������5)�otD�a%���G�)֪�5�PLY������䉺�k���A ^^]���S�}*����g`��ma��	�2*&@oCu���9������X�\\���u���� �Е�K��������'q۟M��[�� �J鈙{`�؞�|�eP�~�!`�{j&$�B>������ 7��*V�|����^�e�1Z	��d@)�B*�
7�z�ܪΙ9
�Y, ����cb�++1"�{�[U��*���P%��Qi�[���7`4��9���<���F���5���똣}K#C�M��v Ͳ&7j���fc༿�l�?]�="��9Ʃw��pjՔ��Rn�,���:+�=o��OmװҹȶM'�Rb��'�)�IZ#ү�6��;�b�蝦;�؁'Qi�Ln���^�n�x�J � )���X�85А�����~{�:�ħvP�*g��>�p�&q�jz�t��Q�r�54���+�3��tY�@)1;mv��ۑ�9���%%�||��})(*~w{%�*ή�}�\l���͏�V||H�����oSY(H��|��M�=��]���z�v���RfP���ņT*�"�qܷ�oqyݶ4:mU��z#������v��~����H(���[Ι����,�[/����;�a��u�*�w�ށ2GC��M�Ӂ�ZY�SPVfm���Yy|�`$;}�����#퐸�p� ��6��/���K��dr�f=���J��8�d0f�v�Fd�:��ߤ�yw�<��Z*���-��<����F���_)�����q�Cߨ��i�g�c �J�p���?I�,E��xc��Ν�"wHRb)�%�DSL�G(��9�h;��B�>����1��$�xxy?~�u�:���T`���ݥo]�i6!�~[�ef���)2$j6�W�����'?�"�����\�6 �q��:�|�Ց?���	�S���J21��ƒm��JpXR-�;|:|�DH��Q	�+��h2�omo��h~��؊��OY�����wL�%q+�E�լ�WM-Ä�o��ڛڡ�G���.��Mϓ��_6Cٞ%nCY}�ȟ'B'��k�s���I���Cy��٘��ʇ�@k�+\�ͳΝ������
LD�R� ��
IQ�M:�{{b���溿z��^HCD�`�]h��ma9�e�E�Zd"��:����Q;$	�?�LW%�PN����'D/�u�ۦ�nf�AY�-u���\#+���b%)!��m�B�k&�!&�o\�b��g!���屍uSȶ�PJ�ׄ�āS{�jj8�P/eT�����<@w	�Zȵ��T�: ��.�z�s)�w/
��h�4HO@m]��%S.�2�s�UUU4�"bF�>{e=at�y�\��Q��~���q4vpy�>��J3!N�������nJ�&���⾾"�.-�c�Q���,e|$�=Wc/�tH��A� �+z��T�W���F�KMG��8s���Jt����2R�<=	��L�#Þ��؆� ��2�f�j�c~��`�{���ze}�j�Bz�v:n��k�}���s�wvv���p����9�WA%Ij.9�y�jl9K�62;*�^z���r�n��pἽ������IQ�X�����x�`#�[?��~�?�2K�s���d����`���ĶY�È���:۞���i/�6|ꋓ����Tj|������×] i �/)@ġ���z�P ƚY]NB���6�H_߽E^Mg����|oHw~� Bh�?1��p!)r���������&<)(#�g�gO�:��M-��^Cv%��m�U�_K�b_�����`A
%�C�X
yx��d1���uﻎ�F�ZY�ߏ��	ԧP�� j�M� �����v��W��A�<CD�ߐ�nl�w�tnsG6[�d�ʹWJ�i�Dx큁�����+�;l��^k4����������
c��d̫uҹ���#�ӑ��_Eo_��4�4H�NMM��ZLXk��/���ļǅ����eϥ��������ݣ#���i���?���~Ki���c���Q�H�㋀O��廪�~\�Ý���^�� <͸ �X�
$xcz*8�%@y�:a}�433#�y, ��p�"���nx�7��Bw��q��so�{�<?=�$�(f�= T��|�ř��������9�&Y�);?wz��?�#����u	�Ə��y�KHo��H��v���V��v�(֯y+8��lhk��~C�f��R��^>��FrQ6u�GM9����8۽������NTT5ZC���A�n�e�8��#Ԑ������!��x�{4
)}�	���R�!s[�Ĭ��0Y,B�rn���;���:��d�v��!cq=��Ǘ(������	j 	Cɕ�u�xvQH�M ��/]���DJ�+���C��e,���� FӘưj>W���n��6l�����G"���Y�T�lr>��4] 8��$�Т�����n�V!2X}s���8<�F3�&�lu�t�u2��@���}Ȇlk7����Ϭ�HCm����0Ʉ��ev2W�*9*ܳPv�Ug*.1�Ŕ.���5y'Hc�FP�gG&�r�=2ĥvg�R6�{�M�V��1Q}��ʢ��B ���͋�ӓ�l֏�]=-��D�"縋�T1��Pl$���C��[�*ZN��6[b��JrsN��>�M��ٵ���{ N�FxTl,k[;y�t�� U���Ⳣ�-ch�Wy'��LP�+_\��ZӤ�c�.%�ܜee��)Ťs�[��9@�f-�^kK$e�6�U?��G��&%`�������D��!��Ʃ�x&ͪq�D�W8��0c�v��f�r�r�Ѥ��~��v��T	;��&t�������Z�Z�e9�f+�49�u��H4���eZ�6j�5�.������Gpt��
oἏ��zB�[�W#roܞ�&��|NNN>�t�:�����J+�Å���۹�e�멹������)7ph��0�-gʴx�g�F���Z��"Q'B�8S�&�|mNC�v��#lrrR��6B�������N���`Շ+����6�L[��i�D�S:ߩR�_�#�4�j2�^���y���{B�@��'��/�kMz q�1t��	�u��竌f ���/���)5_nÊ#ɡ�_6��I����#"����ɸ���J�lƸ�浇��nI�X������{�%Y����K�d�����g�x�&f����.�v(~�e��4%���,�@vT����x��}]@^\����{r"�*N��aww.c":��|6po��}εu��� ([o�u"'��X}r8K�1��<u����~�:�]�|yd��M��g426��1��L�(�\��é���{����Q֝�Q�S��o����s�ٞYc1���@;5 _)S��WGZ �����W7�ϻNo��9��d�=��l]X�R 9�A�@�+�t*�R6#�s�sh:�%
�v#_��@=�ʓ�<^2HR�=HQbAV!�<�>2�S�s�o+��\���냀tC���1�fl.T�풄�hv`,�Ւ5� ]���?��7K�V�~��κxܷ����8�I�K���	LD�]�h]Q��=�-��=��˽���c�s/��KB��C���g���?4
J��c��"�o9vƂX�%�>�ޜ�'�=>������DKC~��A�a�0H4A����l���l���#=Qc1TGn��%���~cV�U^0�i����o��x&ͼ�{� ғ����t�Jғe;9U2����'��,x���	�`J8�xqmAR���NPKr��ײ���h}�Pbp��\�������*dGe9׫�'.����		}7�_0jXĊ��J��g[_7 ҹ��n5^.�͇u�9|A��X}�h�3�+f|]d�D4�ߙ���'��z��om;1���oH���X+��"����;U A+�u�%�����. �$w��-3�5�'(��=H3���^�R*�����
���f�:k�G���/j��d}ʾ�SA���y�����i ݠ�������#� \^]1{f'��Fw@�*N�w�~�KkZ�]w��p���@���C��C�a&>(_�����>7:�d���ȵ�@��^cK����K���,���;	��Y�W��$x�����9�����3o�F�Ԟ0U3�x
���9��&��k���F�2r��}(x��vJ�I@҂|_7�$�Y8��P�N��;�n�C@�n��L�\��m:�@݃�����&��ӓBH�Jr�7�$��l\\A���n�947�Dȧ��܂ܪ�����
FQ]�fEׯ�C�������IE߅i\�o<��*Q� 8��D��R�Ѷ1X�.�>��s��PbtK�[<�FU����@���.ϋO:��F�R�l�� �|�c��9H
�6��r3I�Q��*x� {����.v�jj��"c �����3�q�B����2h���s�n�#��P�!ЃU�FA��[=����[J\2�|+$�J��9{2*L:���B��O���B��KjC;�zρW���	ߓHזp`�>�!�Ѯ2���X泻W����u����R/�����7IO�ȯ��'ޖw��d��}{���G��8�6@��!TĢ��H$�~��S���sBb���l%�BJ�8rWjK��:�Q��pZE�� ��'��Ԏ���m���o��Q�r���ң(Hq@ۧ���%���C���$À���X]�0F0��D9�y�:p*��1��@�F���hq\`�!P1O��*�椠���Sj?��קp��xR]�/��i
�Bk�1�%����rTPV�����ϟ?)K/�Mn���:�>i��4t�!�wQj��O@���1~k��;��Q���y/�����&;3���gLx�!�P=!@�Q�QY.���ZX>�6��:o�N��AƖguH��M�ߠ��p��CyB�@~����Y�_�&�zr��۸'�;�}q舦��zt
�:�@�&1@�?����w���^�H?�!X�Q�p�'�-�+������p&\ �@|�ME�\Ջ0r��Eh���s5D�l����:VV�����Vip/��t��v7�r��y���	Z��74X�/'}��YW%�@r�
��0+��w_l�Z��O]��7a,��bH�$'p㓬��|�j"ݣ�$�7�̋�:�s���xxx &ym.��$$�rP�Gvm;t�9s�'��U�+�{5yNE��� �Tj��c���Pל�*\�1���� ��]>�<�k�t�yxV��k���_��`�����'�ߗvoۏ�|�@��-B��A(@��y����ls��l)�z׼F�[���&�I'����%S����?�A����fB�cBp�4�zF.0�Ho�]��/;:2GM�� ���2�&&���5�9�ʴ�V]�
a�����O}�R<]x���J/��ȴ���G{4J.���<!��;�{gvr�Y�ͱ��W����A'xs_�����Q��/���p#Ĩb%l��m:V��R���u�e���!<�?�&7��~T!S�Svٟ�z��R|P'����A�>�}��ˏؤ'#J��ʔ�K���]WnE8-����.h阾���2W�E-mF�V��Dè��d�rm[��x3#6�#H�X�P����0U{
S���%�f���)�z\J|�@�F��B�2����1z|\h��9N�R*k.- �!�#��a$2����s Y!�G{��2���t�rs�Wεx!x�uO����l�F�<Y�+Qb�m������N(D��춺+�a�y̲�����9j�f/)M�L���-%#)
��A�,)#��O�G�=e|�]ZQV#xB>�ǟP�Z�1���[��������:s#(3�^:� �����h�Ԏ�;�۲U��-�nD���UZ;_s��ŧ0帻�c���=_w�o���<�����sʘ����Oϙ9�Y�؉����K1ضs�>:%��X������d���5��٧�8]������@��8/���K�r<�����WN��y�����>���q����/u�M�JX����#bG���0"�ow�0#	X���c6����Z���,5���n��O�iF�y�@,��iӉ�V�!���w��$c�k��L�3K��c��t�ي�F66����k���|���}G �T��Q��"�7D"+�"�,6 R����U}?��q�����[��oé�l/�hWY@a�p�݇@�<\w�Y�"ԗ��*6���3���7
�;e�ڮb�m��0�7a�o;5NZ/�^�^���h�/À��(��<�8�~���4\��B�Bz\W�н�n9i_�(T�k:��hk״O:E����t=�~�	����	FZ����iNEh'�V;m�_��j�w�
�P^^�z���|���@�:��v�U��v�]ߥ�+Ъ%��b��	{�����9��<����nM<�}~�=�D�%%����e�0�%V�����Nkr[�G|�Y/۞w�B���7�����&�����(�T��8|OR�9��~UmM,C�U^����ol��mn��
V�n�d���*<�
�%J�h�)}��'f��{�� l���D�a��;�#��%7�~�ngj���vv����`������ͼ6%���*���s,$�v���-���ڸ��`|�=Я���o��]�l+�������>7%~�f�a��R�q)nl�����q-}�ef�����m^Œ_�4HP��	���^v]}b���/�[�-JB�"�{r��r]��c���Gf`<Ht뺅B۬\�C7s�B�AF��U����*Ha�cq���ܚ��'���ˍY������/	��U�vO`����x]s�[ܕ�D��r/��KK�9323�ݵ��H���^ƚtЁ� �K�[�9�G-�az�F(��2�/R8au,��g��>��u��n0��5^��	��h��ֳ�GM:��.G��g�й��,�E�~�����U��lSn	UKE$��I\P�g�e���+�s}x1��U��iで+�L�5g4T�n�G}R�ͤ��Ud*�r�~�߁2�����U.��XZ	�z>���Ru� yG�Ą/��#����ؽ�^tad����gi��[��ۍ�(vߕTOl
ؑb8�����ǣ��O�-�ڕ�_9�OGC\�_tB^�o^��_![g�>cvЊvq�7z�gM��J\��Z�AN�=������-.YK�ZV1�G���;w4<��?�9��i��#�bo��	�°g>i��_�-��w2y����t4�@#�'m����H��s�>�E,Y�S�L��K�J��*�c ��D>3T_��***�
��W8�c`2)޳"�@���n��-�Md�������Y1&��̌������g�͖B��;���n��:M�o&�>�sp(�~��@
�����_�z.y�{ Y�X�	�䠲�њ����FY���FՒ;A��#2�J���Mda����5�w7��5�$000�GGR���:��nή�F�?��Qf@�Q;���OU�����{bƱ'�Y��]�|�V���Ό���,��j4	C��?2��*%"$�;s*�a�)�ؗ�G�>��	��e�C\��R�s�=�RI(P�]N�z˽m��_5����D����:�>/�uf?��{BQ�����E-a<�6��>��?�?��u|�9Z����=a_}���}% ��^��>#�f@���%�1�3�rv���QXQ�,$��fe@^�W1{�>5Hcٹ�BT���P!;p�3 �i\�V��"=��P:�3IT#D\\\_**Ї��)Y��D|k_l~[���


Ԑ�����"H]b���e>gp�"P�d3��mF]S�z���Y�U��gE.kNA��+�v����ZV&Α.I�v�(e���BDDMR<e�� �p```�pi��
��o-�o��Ym-/�V" ��:�����X�'�O�J�F����Eb&+����/A&�����**��31)L��CH��w2x�ɩ����v�#��؎ε!�җ%v$�HI,k]h��Ob��� �s��E��S��=R���ԯ7�R����������\�x7�cE_�^E�߾��������y�F��o���
��I0	��6j *�Ϭ��ef#���ׇM[����p�SL�C�2�u�m��>z���#r��c���T�y��29�nb��+H���A��in柞���G�#�*L�`p�LJ�7?���e���UӉ�1Ϟ��R����]c�BY���,	�f㼺`�dm��Ey\ұ����]�gXpQ��E0fX�!�������Mk�8�ƒ|��L8Q�� v�xд�_�?��fQ�3�m���<���LJ�;�|�1��o �~��5���8/v�z���x\������S��O���L翿��������
b*:;A�xd��Ĵ��nU&����!��w����_���4k�M{&��#}��Cs��x'�p��m�Lyfc�=Yȥ�r��.����[��?Gը����6(��n���9H�$g/Z#YZO���Bߙī~.}�� ��h3i^���i b$�7�kW�.��3~~h�n��R�2��z���1�"wH ���{�¾Y��܀�c�CyfbF��&����-��?~��h�n�AؘB:�58�Ywmu56>�7����8���Ň���hw���e�f�)�]�HX@�x��х�T-�V[̨q{c_=5~y����(�?��,�
�I�þ����ܼ�JG�
\��P�S�(z{&�����,;�h��{;−D(U��=���X��(<�ȳ&}f������ܬ�5#��t/�\ssq)<��)N�����tQ�M�zn����w��Ķ�Y޳��6�T��|��4<'ze!�:2�1��`���4{O�X�= ��}��Tk�c�+��?���[��&DO�W�YD�̽�퍸 �/���Ig����`��:�pu�]�����W�U���Q��Ǯ��4��,d� �	砥�9G��4�x�b�H(h��&���$�^(U���F����y�$I�cPkO��S���s���m8�)�C�^*+1 %L��a�!K��EA2�3E�����p��(��2��y"��	Bp+���-�e�EK^Ș3D��cIR�y ��)��1Kԛ�dŷ׼��*��,\��Y��d�49����E	�.��J��0�����\�`  �7]h8�G�+��W;���	�0Z,�4H]�6[��f-�*�2,��ի�/I���ǆI����$D�έ�c�g�,w�^���Akm%�GrE��׊�U6����ճ�v�t������-++�������x���;������{zz8���*;m�1�<P
�a�]@��l��d����%�|Ez��+p����Zy�r}i�H_C��xK�D�(dX?Wt2(�Ea�P�� �=Cɔ6~wM\+��q@��`n��������w�)�A:߁ȇ���t?#`�}����&���]���<�ô�����Z)W7 ��mF�[yO?D�mEE�QD6��)hi�C)��f,]���;�B�%Bw�y?΃
S��Zl�sێ�@�/K����b�P��I�@U�7f�^�>ex;n�Ȕ�!cS��	4�7�B䇺;pm��Fr��d�ٻ<��3؛_!1Ts�ll��̩B�yZ���5��u/O��ڢ6�*��1��GIRbNyM8/��p����\tLAL����5�~�3�H��ԃY�����z���q�t��)�����+��4�������]���䤖F�o¤K\7�0��43錪��K� ?�B �μ��_�1�?h!�^˶�6��
��.&�����F��Y�ʖ/}o� 	��;��������0��!�()�L׻�߁@t��r��)f��&��ֆMq
�ǻ������so�̂�an(#�������	9)��n��Su�����^k�N��$��'��z�j�S�4u�g\���H��	,�0��HMB���GH9d�j�g�,���ת�3/�1�_�mk�wʼ`�C�TGLC;b����� ��{W��ug��C>��6s���x&۷�Z���ON������"/�1��κn9��%;��5��z|�>%d��XHaI)���6��Yj��������15���Q-@\��J�5X1:x�������L�FAii)����f��~��U�(�9�{��8"%N$;��ѢM:ǽ��9%$�
�3P���UR����_!ߝ"h,�s�4<�d����t����~�����%��%�|��_Q�:��D.���	��:.9v_�_Js��
TF�~�ؠv��L�P�"_D�pjV�0��|H,��Cڜ͎��z�������q���� ?�!�������k��KW8p�ox-W�֦7�{;�8d"G΄�2f��|�k_�Q�毬�o�)�$$\�fnE�ԙ��k�YW���)Z1�k�p�����ي9	�|F\��N�u��*K����ܶ��~�؇��7���h`�	W��ӑ����P�yPq�UFA�->�+C<��u'��ۈG��*V���S2&%��ɚ�NZʆ̉�s�*�����Y�U�L3�����L��_�K���l�0�=��/c�}��˘x���@��ڎ�K��{n/���ᯪ���B6H�'A,�����BA��ߔ�o��r���p���p���śY�,5vΨ��㤘8;;9	�{ �G_Yq?0SH~�t�����L���i�l-�Z��[q@��C�Y9:t�~ӽ�4��М�ן|����ʙ�����/0�u¿����I�J����5$N��p��H A,���A��ɓ6�E�����L�hЦ6��H.��h�ėH�T�arq1ryYhwL�,�"n�R�S�M&с��b8Li��QD��Ks��9�q6��SN�uB˂@��'��5�x�F���6�J,�fc��O1���K$Ss"~0mN��,��5�a4�i�&}��ᦦr.�/Ӿa��i@�g,���yBB#�4[Q(�:�CI>��:�S �G�ӡ$]����F�4�P
�5�蛿�ǉ?|��Jq^���W=�Y�8��"LJ��x���l_�5�2ב�3��z�	!+۱rX�fx����"Q�趸9��[�Z�*�P��ͨx��Ge�PX ���,F�?����3�%R��@º��Y�<#�ka�̴��Vx�V7���;���'��������zV.pA�T��[a�&�5y%�P�la?�pF-V-�����(��	Ϙ�d��e� #Bo=<�:��Gj�����W5tXSH�]m���Ts5�J���}�ރNA���#$b0!���?����g�:ʓ�<=���"7#z�`{K3:ԡ�#�=FS��� 2[5�N�4�.w̅S�q� 0��O��'o�k���:��T�/�9@������5b�n�&@�:��9r��^�:����PPۇ+t��
�y�_�@�:-���m�ZA,�;�5=��+�W)LjB��5&3�X^���w�j�:�l��
�Y-ܝ�����4I��9��-x*+I��B�q���DA��O�?%e�^��v'�a$@v/]�;,�ʯ�J�o�(0�ʃ��5�	��T�����@	ǌcw#��hR���H"W�X,�a����[��Is-�ƊȜ2���Qi�Nv�Ci�W8`�L.V�J�a��	Jvɏ��C޶����f�M�qȫ�,tf��=f��F*�E*Ѩ��������'fgC���[�$}}Eb�.^!�.`E���b�3g�����ˤe$���e��4���S���#�_��"�	[D�NGZ�.�d�Q�H�Y�%�)NNN^bW����뙦���@��H׊s ��.��e��]��!]�j�������OF�Rz��i��$���ϭx����J?�VD���Q�=���W��%� �!��!��1��-��())�t��]A&��IW��3�K�:(<�R���Q��_�_�Uv�~� ��d���Qv{��)N,�{��3Ƶ�u�Z�a���'�k�Zr�z�x+�k����?�o{Q�����Pt03BܘR^���y��cJ�i���H��s��� ?�=�oo,	�aM�oZ��K�v@X��(���e�ۊ;����tk렐Z�9x��C&oVH��#�2�Uيc{Ӌd�*�	��o��|ᠣ�z1�Z 3���>��#Fra*^WK�?+���w���� �)�S4p�vZ�۔q�᚞GԒ��Gܿ�����_�P����l�x-���=Q��	���e��Q��B� (��B�K4Ѫ���'�3��-ݳ����r��(i|��,�|f¨����������B!}���&��!��ϴ�.���	h�3�W���d�d�d��d��@Sww%���CI6�`?Ml�	�K��2�ߛ0���Ɋ�Y�X��.T��)/���eP��#<��1��2��!�W �Z�t��÷T�z��%g��bZkE�o$>7��������)_�Ǒ�+�O;�1^�tZ���[�
��N1�9U~
�B�0>�<�7Wd �'n4 l������@�4Ux�l�p>���x�H�������P�%���%|�,�5 ��Wc��+*W��>�����bF�>����}�rcK�׭w9Z0{�����H&y�7�-�V�p��pc��m�x8�jy\ޝ��w�d8��L.�s,Ч�~�@h^��4lϕ�a'LP�ճ�}sF��q�5��"�,��c6YR�z��fnja�r%=(3l��B�n�9JVe�q�)�J���m��C�ۦD���쌏��'Y����^ /���u����f]Q��-�+��1J� A��x���?财���1��d��rI���_� �ʹ\��\c��&��8䌬w�G���~���WQ�r������ ��Y-�2 >·��U�*%?���X���P�a��(�/N���&Z��Ac���Y��PEU�R���Oo��T�µ{w*$+�J~� nv�F��Ψ�+D�`�A�	�G�n�)�UQ�ht~˅9�䀋
�t��I���1K՚`�!�`'� Q$���Ϟ�#����<s�[`c�'�Op�&i�	bø��(��(~�VS�X�O��b"�0�%M�K^��ʴ��S��U�>a^_g[В�/��6��D�- ��x�l93�����PA�9l�+)>��z���`����g����[�k
�~օ��S�Cb_�����7"YPF���kcb�h��0[<P�嬉�n'��8����;�/d�c����b�z�NP��ޅ-)�r	��I0��xi����xX��r�s��>m�����ε�$�DD��"�E-J�����;�Q��D�]�6J�ha�т轎6�#������>����{���k���Ȅ{�g5�SÚK|����y�'�no/�遳&J@��*_�:���1�9�v!$_@�����!�J�d@LQ֋�w���� U�i(��r�lx�M��U��p����)�%d��V>���K� �O�;>8�TC��b��\��$��9�������7xy�c��"Q��d5��s��~�A��-N��LN�d �IR���@�NS�'��������ׅ��l���Y_� �?lB��yw�^�2'*5�(�Ց��-����ng~�`��`�p �T�� D�-�,a��"�Rs̉�IV>h��6����*�����!w�[���bx�a�����}r�{z8I�$����
 Ʒ�Va����o�����ϯ�k�䳉ט.f5��9���, !���A ��!�	Oʇ��ĸ;�x�C�h�z	m�]��5܅�G$�� �=ȁ`K�Gu$^6���S�R�Y�E�Y����Kc�����I�t5���L7"�s/�W4r�?P��3�`�qO�f �;�C�?����e�P qH�>ݤ:%���ѷJ>q-}.}�M�j&��r��[�+�-�y1��Q���O/r����L,�|?���
U�;R����q�Μ={0(i��t`t���ߐS&���&���ۍs�oO~�"�� 
A"̀��w������\^G<K�y!�\6� ���&���>8I�~L 兵"�XU�h3A��<��@U����ZV���H0\6��Fdʛ�Sz���񄫣ף�S��9'2�W�^Ú�r�ԥ��u5K_��Z&,�-��������M?�}���?m�S���Y�<%�9����vRki�g�Yw��|Ի��%'!Clxn��~�m0�A
Plp���%�˰}��D�
��oV�Q��H��ER��Ҵu��
��K����{�
�r���%$�]ox� ��\$C�P���1�,�,�R�q��@#h����O�237D�"k?> n�9�x�PXwT��¥��%�����I����~�[�3�q��6%1p~4�[��":1H�K�cL�|,5D&��T8��^G�*�ǟ߈�l���]~.�b��p d��/��w��E���2�|_e�Ȝ�V\�d�`�����g��'0	��Ck
se�j���7���,ֿ�o'*F��W�P�WHѱ̑�޸殭f��N�.�+���H�>��h�s%F�u�	��_�d��+H��?A��^ה! rZ��,�2�(�~��ǿ�3cus��o�T�Ix{��$��r���^+����p��#����呡�1J:��;�\\�H[�{��ب�z��
�ai���%<K|x����7D�㼚���Yo���#�)��U��:�>�ר�򏁐�zd5DV�#�)s��}3���+b�~Ne�35��)�������v��zg����Y��1]�k�{�)���mB5f~|���&��T���#IL�X�mH��l��OV�8bCD��3;����Gt���<�T}���{���yg{�Ckts�~��P�%o��ǎPV����	�%xG�s��NAI�i�e_R��!��4�)Y,v~<k!,��1��ah�ښ��a��ge��������)� ��d�~T �H[����WĹ�SƯ
 b,k���BDpӕh��.鋵�Zkx�C�ޚ`r!L��m����q��ǶFr��^"D[�⌸2x�%WnH~l������Y��{�\��o�J����G�ZJ��\�gɅ<~������UU�h8+.T����}�H(�� "�$�L�n������r�9��+Sׅ�`��Ef)��׭-������>%do��@�x�Fm�s�������/��vnY}�	G�R��pi�r䘂�s��{��g�����?�7�j@�<l�ueN��\w
�������uV���m��a��k�����D�K���&�i�s:�mp�m�A$�T#h����Џ�7���À/��p�&V(U�2� =F|o< uH!�IQ�����k�W�xs����A����=dD>^�,���`�P)J,�}�I�^Gۈ%��	(~Sɞ��0ᴑQCԝƀ8�p�/�tNǖ�����[Kx�:��9�Β�+���u^Ѫ��El�Lq�A��w��`��<�
�,U�8%T�c�8����ӘG�+����%�jM�L�;���t�6���3�---M�U;�u��EyMO9@��v��i�L���������,U臢c�	yI�1�T�����¼��l� R%|�4�4��һ�	R�,|��ܼ�H48��a�����DȬ��vi&���z!�_*R��~�:��H�5�I���0�aJ�	�rΩ�n����h�����y���u�\�Z�D%0�6د�US*0H:�!���4�fn�Cv�����'<�=�L�r̀6V1��uYh�����X�� ґl�Rm��B)�l���q��<���įN̨�V�����|Gl�黀zp=w�u��n��+[�^UO�uIV�U�qR��o+J��O�P��e��y��c�y�l��τ[�Ʋ a��Cϭ�=��e��z.�����ZN��GN�u�o��Nd�ʋ�Su��U\�����U���� ��^ ��ஆff�<�� ��K�UB�/bw5Oϫ�u�$KA�g	�w�TR��`6a�+}���V9r_���
��S$x�;�����ؼ8���8Ċf���$�)7DH�m������.Y6�񽧱LŖ�{�����Q�zW�Uz���0��I���ҹ����i��n�'�DT��c>GIj֓�W��'@J�k�iĉLjp�(���yo���C~�/��H)qh�bp˲���q����L�	Li��U�n�_a��F@��M$���9�"x��S�|o���iL8/���Oۉ�r&�t�L{�)ӕS�m?a�'̃��-�𰗧�Bh2A;R���k0���:����VN��g�U��B�R�+7l����V8����x�p��lf�h?�o�Xv}��B��M,Տ6h�$Wg�}+W�P�~��yˉ��vPK��G��[�����K��X�����Qp�����g����H�޵�#��a+gF�����X��jݙ�C8���ӒZ%Ͷ��;/���U�j6��9$Y�4،<xv��;S�0}�iW7Z�A�𓄈���?�KZ���7����kң��B6���z ��$S�xE�U!�3��w�8����<»l�	{��5g~���[%�����ؠt�e��G�b��&Y�+�Q	/6q���66�7v^-m��V�ӿp����n�x$��ѕ0�ל*�HT���g>�I`J$E�����un�x\�n�BK����cޮ��PH�����Z�f�v�.���=�UP��'bA�48p;?�I<5�-Nт�ͷ���j��������$kg�?�Yo
�yn�W8�g�l<�#�k�K]
jrn�)�����������bq,X*,D���ZYi���Pz�4(6��]��I
����b.���{Q���E�*��]�����+��{�/4ǡ,��>'+6)�N�S6�y,�}a܎8�v��b������ /{�8�p��$4��w�*�g�i�]�f!u�d=qi��on��wMI垝�"9���$�~vg��[�G�m3�k�#�$H��]�=>O�T�^���8r��j�T�&z�zϫa�cz��:�ƚжݧ0�9�!E�VǢ�"�Pwا�_%�KI�#���X�ٿ����r4��hߑp��5|�3(s�N�����e���[��+��dL�:�3�\�?E�����	,�J�D�Ӡ@�QK�x����WH�^x�6jإj����G�v�����E�b8N�OX�3�(�q��2��D�K_��pvRjE�d�jQ{_T�74�E�k?|�ΒG ��7��ݵ����DG��I���H�S>�+0��R$�D�����d��gg�j�ƊUh�S1��<�z +�&�����D�=�֢0�_������o��U?ܚ�D�S-���L����d�` >���/�Y�abM��p���C��c������x*}#B�~���Ձ'���\�+(t����5��������P�S#���3��(��
j�Z�D�9V������ޑx)s8m�������
�������`�7�Ӣ:�b�۲�[��{#[�i߮,i�iʬ�^_�%Я7�3 ��!��B��UoYU3�*���,�y;�Ǉ���k?��~~����{r����	��w;K�vC�����fp��Ș��E�¥�$X��)h>vb����A��E�l�ES0E�7X��˹�O#�D�����I_zH�I�7�R��MS�y����yv����B��v4-0"IZ�5{���4z��2>DN�ϯ��O�z�f�G�~�=�:>�:�F{�^}|D�sr��w�#W��)n0��Z1�E�}��@L&��4nc^7����y�<�Ȧ{��B� !�(F��H���Z��"�K�9��.7ݽx4Sg��\�`N�ϵ ������ՄƁ~g���C/��WS �X�_+ڶ���%&��ү,t�7��p��%� ��Z
�ri�~�|B*"��rP�Rq��R4j#�1f{w��W��J��~5f]C��k��r.~�3��2��z�Z��?����3�3�m�.��Ȱ���C����,T�o�#y�2��@��Iʺ�,����j�Ӡ�g(*��l�D&/<F���H�e����|(��3�;�{�gY����]���n����{v�T��~��k��հ�!�!��t�(3vA�;�>��H�s�=�q�2��a��Ej%�j�ޞ/ J�����{H�5q�r����;��X����d^�霷?�e�}	T��x펬LtZ+%�i#���0�D+ekN�e!/���EL�n��,^���4H�'�J������F�����M`��yw�Κh)tG4p����(+#*��E��J����E֭*��b"m�Fѹ����h�JzI���	4mԝ����� �>>�t��i�T�&��*��KbS`�r~����v��p�⅟kv�Y$�m��#�m�ݟlm������9{~�����R�����1ϻ�;-�̓�	�ͻ��F�,_�K��_��;�fm_�.�f�|?0���T����(/'�d��|��3� �~/,�k^���	K�����}\`~ZS\�Z�~���K�iu�~�ӏ)�%#}س�` c��@*�0�K۳�5Y��2�Kj��0th������$QV+uUuW�ũ6��)���1�r�}·~�뇤�/z�'�c�	s/~wȔ�*!@6���C��n5���O3���y�8�ծy�ó���X^^nL�
HqV�b�F@��x�jKK�!s	��'�������g�����6q3����O�|�/�d�G�ttt���(���ٍMf�&0ڣj5�j��d��ϹvO�{�i�C����Med,e���©II��Un�=���]2���nԽ�p��l��g�/Y17IF&��IePx�g QW&�;�����'�a� K�>�F/g���@��~<�Ho�?l f���G|+�$66��U�G�Z��
�9�e/�vo�ud�61�_W�<�ݭ]Q�눿PTzz��B�F��IH��P�r�Su�����t��?�F�Ww�t�U0��SB��tl�gW��+�IC���qE˹�LX5@R��A!j��{B�"ڥ{�n!$��%~Y�F!$�~��x���-mp9w��s����8��@;pQB���|S<����G&��e��avE�;�iJ�gĺ`�H��W�۳�r��ץ���I��}���ˏ	�i�� v��`YX�B_�4,���,Vg	7	W'kMp��#`�<|wiip+'ArX`_eD�ش�W�vM)G�+;J0O�}�.�`��|vDr�U6�����(Fmf�ͩi@��#�vK5{��*n܀ԑQB�L�pwo,�E��1G�f,9�[�}���)�M��4oɿ�.��O��s�w�C��K�ل�"��f��$&�s�{��*L�e.:�𘅼��7u���BS����U�Z�8x�4�Bmv�0��;ڀ���#�6�����ￆf/���7� �x�[  �t-o@�cq���U�q�d�8��]���< @u����k��n�$�_ Üs�Û��r�������+攝_���eb�k"�/�MP_.��]#������H匓��S2�����}I[[�{������T���`/��H+0ᵅ���;�S�E&;�J�5��U!�9%A3lh Z����:-&1[�T����[hH�ܜ(��^� ���y3d'ʔY���N��=�	B%n��(��!�Z9��t�m��j�$|)�/�L�7�B��źz����=%W$$����2�@�>�M$�Rd���Y$�rJu�x堖��+#�49��Fj�z��y�l��= X)���^��"���OY��%�SpBm^�o�j�������+�е��\^���E���t��W�8�fu%��=�Ԉ��S�l��l�Ŏu��2�K�%�	<y�|��I���?�q���RVh�Ӻ�+��w��2�dHh��E������\*I���S�ܒ��C�ڞv`K��t�H�H��A�E+�Zos��������S�<[����nW��t��Zp� �z}���}Q,�(ϗ ֩ۄ���(�3R�_�eOn�4�?�TQ愠�_N"x�L�Hu��J9��YH*ć}S�dp�����3�O6� ��`�p�h`p]BjY�P���t�O��xI��I��'����y���]��E�:��VNo7�2�%=qu���.��B������	a(��W�#�̊��@�Q�����(�e9ۡ�yQ��h'�@�\�`ޝ����s&ƚ�@��W7t�!��ק�r�A���]�%�nPJ���S���hK4���1�/��y3X��,�I[����Vcq�mq�Qc�ת���NVv����J�S�~�-��H���T�a�A�a�^��j̜D��Gb�\�+�����%3Ͷ˫�y����RfN�:7��#֤��9'���x���ɣ]������̸�|OiCO�,�y�h7Ck����#s��sr�$K�]~�:�_��~}��� �Rvf���g������i��l����v׹��Z�Oq��+�v޾OW%Ѽ�z���W���wL��a9�Zws�Y��W�����K���f���#Q��#��+o> c�S��)r�ۮN��pb��h&It��$���ؿ"��=:jkBK�K\�[g��z��^�&�mP�K�H�sB�d&v�<��m�v8��t(@���'S�8���L ���:��*���H�Tڒ��+-�9qp�͹�V��$=Z�I�,��|�<���t Q���p�_��J���ěK�6B� �EE�>�lki�#��kfp�V?������ߴ�)��_��u�s|*!�uj p�#���/��B�	�g��)��n�P��ig�3������������R��@'A�FGt,�@T�@Wi�	D�\�E8���hF|���x�������g�s
��F�s��ue�j�.�5ִ֞��܃��&�V����/ �J_��6�)⟬��\}G�?���8k�!���)O�@��[W�RJH����m`E����ޠL�ߊ-��	��uR�ɜ�¢����3��ka�\NB�ݿ9�ɞv[�!�D� �{�R��ǻ>�5Q�.��s���|����!�<��;�_�#��l�9���� x�	��zmd�ڨ�ċ��+|(��c�)�12��"ӗ ���%���uL4.�9@�@�>�=�O��M;�d��V�zz��k��z6��=��"���Sj�O�����Y���c;�	��J�R���OLpМȈ�- �o����5��=xo���cN�2��{��"�ӱ�p�ٚ����|y��7u��w�){S�SHvx�L�<����4I�h��)����U'�ojH�kd�?*�Y}�� �h�i�ƿ�{g�ÅM<���;�=�8� 5�!^��}�a�$L����': �%�&�S����f�u���9��C�9G/r��{H	S��^���쑩+M���Ja�/�^�yr��nOXܫ�4\�H\��ϯ�Yð�)�<���L��O��<�~���!��?�h��^D�zs����N���kt�}�9,O�";�dL��2�#jt�܋�;jXd�a!�|����sCD���M�*A��N�}�|�`���_/�"a�»�e�0����v�Bc��Tc����M$�g������WA2�ą��/�q	��)L]�P�p�J)
�e�y�^�g�^�?����ZY�f�,��i��������܆��zٳe%��������_�� �M�;)O�a��1G<�f��>I"� Eל܂��ã�g��Y�j/�S�wW�u�7�t�H����ιlT�-n8J)�?|]��}T�}/�ѥҸ�Fä��¸a"�0�˶)��9rɹ-����<>�~)�3�K��礑T\S�+�����]��"�(v�P��^#iJ"�$"30GK~2k;�5]&	����*Yu���^F�����d^T���|��H�ۧV��=oO��Q��XI`)�k:��V�G����Y6�.�Pe`�Zd�ZId�ꘅI���U���8�_RR�1"�;N����!��b�nI�{��x�=�L��������0{ִ�ɧ'=�������2V�,���?,]��0����\9�Fam��q�?ZfnP��c��CT�qY�5Zߤ=}�7�q\?n<��A/=+2��x԰^ �������}b�Lf�U���*�Bv�L);�Z�Y�5�ji�p;^�	,��N������(��C"��z9�B%z�mu���,,��\���q�>�3WqU��2�������j~2�YLQO�n�L�̆����"J����J�\6�AB85Mq:σ6Mc�J��+˜w������5��TU��،����!�������m���gfh��[D5��@N�~�1�#�ןD��o���Dw!Bs%d�s,a+�����h��@	��Eœ(���r�R�7�>�T���#��:�A*t��fr�Q�*��ścFUa�͹��)��vm���!f��̥=�ʽ�Yy�
"��\'`��NI";��~�e����v�c�0���#���Пw�~����8��,- /u�$]����؈�&�I)N�1�̪vЭ�U\ Qҗ3�(=�hկ��(d�t	���o�S5�z)�r���R�R"D=[�ۭ˽�^���3�4	I4�MÔ��y����W'���^.hfg��;���s�����k�y;�z�b�/<���'_�
 X$��wL��\d�W�y� ܤ�C�A<�^�Ɵ�s�]U�@�N/��s��5&�D���Q�J�Ә�.ȑ��:{^~������F� DeM��n-�9���r�����o%`����Y��I�9�w�|��5-�$�**�E�4?U��ib-B�����o2��-�e���<8��z�� ���7���d���K���&�Ԃ'c��b�bF�A�jA�\�M���5j�q�1=��K阨F/S��y֎Sh٠Ҫ���xǨ��Ev���f��r#���&"������i�YQD����o��W4����L��,�#�(�־)|���&!yR��9�z��x��n���co��Q��sEc�I����Nc��8N3�������)����j�n���R��8WcE��#\s����b̬}�e�b��v�Nz�.V�91m�� �qֻ�r�����WZ�<?ڲ+.��E�FbC���Q��JC���۫/�V?>+�����z���ʶ�&1���nfNm_֜����-�԰�sLm�M�SL녚�if8�vFUŵ���k�k~{*�b֖���E����� LJ.Nz*0Pf\^&�����t��ɖ�;=�M���Դc�'�8����5���YF��f�~s[���O����;'�7�53fǌD���zy��=I��ζ(��F�e�Ȏ�=��w�E_1��K���l�>`3�c��'?���1�ǯ��(�ְu6��A#��K�o'�f0aP�3�� ���f곁����0mH}h|{S��A��ݒ�[�9/�����P��G�Pr�����+�/O�o���E�{�!D��������q�
�~-M��s]p��c�N��_��9��8�������g�^-��}3��;X��˷[!
�7_nEas����]d_cs�8�-[�Q/׬����i�
�Pފ
~�,�Ҧ��iD4�4C/b�O~��R����L���I�^���e85���|�QCm���k�������,�k��J���]@.Cx6� ��72��Wrɽi���=4�m�������37�r\��4��dlf*4f�i_$�F0��VO��N��pY�m�F��H���e��*�)&�E���ٗ/��o,G�M9�T(|��YR/�5��O.J�eg�Qy��=��`�"�L*��v�[��WW�F��)}�����#��tJ��.�5f���"����	����K^�)�ń�Y�e�E[����a�vJ�4_���~]�h����"�>ן�sJ�X���.�^����s~&�b%�;
6�I c��<������%�nS.u&@�e�z����P���p�H*�45(�'���=��KґU/oU���}+ KʮpF�7�����Y����.rܦ�%�E���gL?#(Z��7�����=�6w����ȝ�\y�3D���7�~)��9z�6�^���S�Y��ձ*0#x��.w���F������Nl6�w��|�����Gis���3K��$���J�W��us�x!��L����F�f��,WGz�J{3�?�������?��6�D�%�� ��v�n��	��d,�X�~5L��Tvz=5��t7�����TE��nm/�x�vc���y��l����5?���:=b�F״��5�X*R�k�9q:\�]j�q�U���5]����T-�&<�r��ާ�!�4.IH 3|Q���\�.���]�]�#��Lc����� '����\ը�3#\�����^�P���&ڭ(A��5�/�I��jz���w{ZI�u��ȉw��I��5j�W�l��^���3 �ȑ3ӈx��:g����G���&����/�وE��D��: �:�R��M�e�FR�_�Q�7��\�����zp�H9��C�ҥ�I(-y��kg��Y3�C$�de���IL���'�C�� Z�_�N��&���XH�s�D��xD��z���a�$;��Y��������ҽ�5���䏻�Q�l��PhZͷ�iu�����Rì϶i �|�NW�T"1>����ƾS��%�#j+�Qkd��U�`�ข��t�۪��('�W����̰Im�ġ�`�U��J-��D>�l��%+��O��8zE��u����E���`l#�>�6W����fTȣ'���ʔ=�N�'Չ�� Sm�sf��]t��b��\a����T�#�2�{��Ib��)D�JZRȚh*�z�a7�BWf�x	��
+�z���r�}�A�gN��)zѺ��f�ڴ�`�FD�?V��[�\�a8\���g(��yS��--�h��26rr�������(��������Ym�ѳ*e�dv��h[��I{ɨ������\	/rŸ�z��u��'^��t���J��4,ٿx��5W�6A�:��&�*�`�[Q��4%��ڿD״{�[MT���"t�,�*�+b���A��jWP�ӕ5�!��>�H�J{�~
S�h�3Y�.F�$5T�57ؿ�gD�˭��F�5���Z�tu̎�=��$���j��E�CL�N���ᘰt��.�F0�f�g�5��>f�c���Z2;��*г�Xu�\��o[�7�q�Q�6c�œ.����K�]��_�]
�;6�Y��,j�ڕ�]���=�@��6z� �v��k�x�����3�o��nV���e�k�w�l�B�N�F(`��Ŕ�j55%̗L��<ཹ#�ͥ��H"���;ﲬ79ӯn#�J��4<g����ɰ�,�z&ŝ�-���U����Tz�&���3�x~ś�����)z�_�HC�5W����OEO�^*�z���X>��*%���Uva!⺿$��2�b )���"l0�e%��̻���7c�F�/���:{y��O��gE��>�|"��6-��L:)=��뻁^Wv�{���%+�o_���{���!5mb��h��l��bK�9��	3|�el�ky�Z��b�$BV2o	�[y��jD�(��ѻME���W?���k������˻ޛQ���D�FŠj�߱��w�/�w�0)��i�gP����=	�tK�iιH[�M$�JP%6�a����|�K�sK�\�A������H��AԬ�V�ط��O� �-?;���R��5b�ܣ�/(����T6�)ϟ�=Ғ'j�*�s��zM-�*\�?�-:�k[�{��j������3>����4X�^q5�7z��:�l���T+��3����d2\��5�B&�jW[|�Kz+\{smez�2��$��X7��KZ(�����/v[���h��l��q-��k����}�E��������`f�`N��A����\�ppWRe+HM"AC�΋e"��@Frv7w����n��f�?E��Md��3�^��^|�n��:��=���=�]�2J\Z�P2���~q ����Y�׽T�sƪD�f�!����HR�D�URۋ3BZM�4�u��c�mJ��������r.�34�)���[R�~���(ql�2 \�jGӬ�85������;kV�Fg�wJ�߷��G�f��:��^YU����i��k��tB��5֨%`ֺ(N�?�.߶v��/���-;��rev=�jp�ތK}<5�×7Q�8(%�um���[1��=�E�1E��O��_β�,~�?�!(��
��O��eS����^V}��l�-Ϥ���Q\�+&���tGj~�xn�g�� o��̟�ǓsGL�ڰ�0m���_t�&�K���,��A�gxw����N��+V�/fVx����Un�ēY��-[tDzv=�{ Y�W��}��Fbɯ-�5��I��<ǧ�"����e�����R����7�?��7�{c�E#��K�$���D�{˷�G>2�6�C�*�ij�p�-�]��Xad�C��c�?$QGY�(s<�����ˈO�'�d���X����q�U�����S|D�����8�mI:cQY��̼�BM��ب��o�g_Ҭ����-}pۛ�+���|p���*37�.�:�Ƈ���$8ު8�B��X��9�>���|�t�#*�s'�m���ճ%�Y�lr�� Ɯ��3{C�O���֩F������6�4hح{\uHW5�=R�i�����m���g%m$��~�R��s���C���~Q���
�4��n�R�G����L�	*_�."N�M-��V�s����p�U�	��;�b�J�xp
�ZUe�j�}f�/wN?��5���#+�:j�rx~�=��YU��_:$Y�)�8��*�£�@X�����1I�*>���<�w[-�jn&N|a�s�I?M�_��Y/�d�j��3SX64u�����!�燜}eM���^�U��qB&���8�x��V�����3,�Դ͉�M	b���%���xGe���^��ON�MiZͭkb�$�q4�\yFs
��N/�du��� �
8��M�L�q8�X�����zH��3���R��z��e7M�Q��3�Zj����׍���Q�@Rb#���~��ٓ��[[�OZE�³��}OϞ���G.D��kZ�<(���"ݐ,f���4 ��b3I��Em��x��2��I�D��U?m��Y<����x�nizp����*��ob6'h�'��^��I�I寊�i��=�qXX�ĠA;�U�e�\6HL�+������--ĥh��gL�^P§�fc$�S�6V!��?���(�<T���OYz	��Ϡ���t ��j,�����	]����y�)�3T���f��dJ�Ta��vH��GQK��Jn]��FL���".��(�;���׃�y��j���n4Fh�]�_Ӳ�����x����Z�ɪ�^�rv�����`:;v�q�||���˲�H�ll�<��Hnï��]7���͚9_٫P_�89���yZc��M��gԡ�l�>����B��:I��݉�'f�7W{��M��bʿ�L�ge4�G`O+߿�q�Q �����r����/o��"_p�"�&���&�4�S�>k�*��ϔ��MC���5�N0	��Y��Ь[����O�3J,�K6�n��;�������5��DT ������=S��d���p�B�Q�c�S�_��G�ElA�|���b'��e���M���'5zΉ	�&M���ZG�IG����,�ɟ����Z�G"�b~���w�)�,XO���5p���X`�%7�R����+'��VY�P��%���cSCַ'Z�8�l�;�g���!�5.�Va���Qm��<Y��<��،>C��}vA��CC{x��*� �e�� l����������Z�ʆ�	fW��(��}jEE�ZT\;GN���ݻl�
��맷� ��G�����,F1��`V��
s3�� ����s&�F��^<W��&S�$M�dw�?y����������oZ�5��n� H<�L�����G-�l�<�zU��N�ȟϝ�}�ܿ
N�h�8��� �#�K(�^�����N��Ls��D#������8���iN4�$n8E#���R���Y��Uř���U_�4�q>��_ZJ��H�r��J��i圭��iD�S͑�5FJ/֩�+%�D�O�d{�{Nώi�9&E�F�E��Rc�xn�
;1cc�	�m�i<,ad?�h@�	��r���S���Q�}��ȟ�;�����X���3/]�RVFƲ�&��^�gŶ�iw&��0ă�G�-��z��Yۭ���\�SqW�{�߄����G��L�j-�l���UL���>���N�%X\��`��;ZyF��ŌV�:�y���q��pW�?�x��u��h��`��Q.�?�����	r�`{D�^vf����*�E�Y�k7��#�!��.kˀp{����ʧL�~m���,$����ZW$�9�h(�>&N��;��6^U%٣�N���%���-�~�u�Y���$�=���� ��"�����`�'�G�C���>���f.
S��N�x��$b�(�޵�ļ��fMڣ}C�=9}:�v,�O�����ƃGO���̠�)�#�ç�f+J*�b��F�"uJԮ_	}��nj�uV#���]%�.E���@�53X�9�Z�xi����n�@�ѱ[���Qc76��9��*�@��*]\�'84�r`�K��Ց]v�~�lA|ư�־˜Ub�
E(ILnN�_s�����Ƣ����Pm��D5h�E��ޮ�V��i���M�Y���jɇ�zi�<X�w���f?����z����vc�anf�^< h6��ϰ|_�V��3�k�r�(Y�ҋ�J W��?���Eg�O���(a��
dH�#_S��
fý�"ECbHՁN�:��AVL��L#�v��p�Xw�t���֚̊b+ܣ=�31�\�����KϮ�M"�|'�h�g����Ivw�0qԩ%��G}(Z�6#�:��-�q��y0�0��O��_���{~�_��F5�6� �m�^��+Z����3\��lO�� ^��g�t�\��j�dİ��b{�N� �QB&Q�ܿ�I��lS�IP��y��	���^G�����k��D�=v]o�-�c��G[L�ݨ�A����Eb�Sv��؜�GE6���½�����y�;;g;� 4�wE�z�Xy-1-�Eu4�~(�Q��`zl�'-�
X���4��`+�)����<�+�H&�i��4�x�����Q���d^���va�Ƣ^���5ܨq��H#O�)��������#�uPb�xH}h��"g�w��H��Ѡx+�)m�� ��y���5$�l���?~y���frdDo���2^Ջ*3D�S�0 �k0����KK�'? {��Ta���"�Ǻ�"��8��ou�h�!X���+P��O@���&�[�}�;{_S\lD�l>:_��
�3>Ϳ�|r��"�8�le�1{j#0I� �4�k���M�����v ��º,�.�9j���նf;5�`���d�l �2��w����K��mYO������/T>�!�"#���Z�����I
���O^?R��;Rq	��z���mr���7[�ۀ%��?��ߺ�0�V�b��9��6�J#��pZv6�G?����C�`�3ZrPAٻ��I��$Z�#M"<w�-��f(]�����C��0!z�n^�Y��gg�Tc�h�#��E'�������Bn#���I���x4^�(��Nڻ�z[�h��^C�Wo�$X
�����T�}Yv���*t]ݽM����_J��.9*����������eVf�2NY �/<���p�}׷j9��3CӐ�N��9�ɻ�,�0����iX���O�F�ڿ����)��>팆�~f_ 	dSn�:ܪd`vXf�x�%�\!�>�B"�0�����A�R����;1�H�Q�k���cTORB�z��̷L��^nv�ަx>��5'�0u�Ā��lBW�,�
����<�m&�:Q�`��M��g��u힧L:5X=v���ƯN���a���lA���x�w@ߞ�9��:��A�"	��r�X�S�Y1ZaU��zq+4��6(��݋������fA�\�3�Y��.�ftl4��MGpQ>��>h��:�ԘV�k_���׾��C���ON��)�hEʚ]�e���e0�!���,-�P��c��+2�c����c섌e��۩��\����s]���]�羟�r��L&`NZa,���6�յ�?��N���b�����8B{�����(�}�����N�E��uog]�Vd�����%��>ĭwBw_�G���އ��UT��h�Wu���M��D�1��Mj�V���Oy��sێ�3���,�^e33�l�IT��I�|�����/<Q�N}\FOr^ttc�&�������w�Un�G%�%M�m���ѧO����+1�O��"�w񽮮�K���a��U-�+�k�����$�Z.�tT���+�ZAs�`���G1��l9KӰ�hc�W����*���>��b{��2Bi�4|��!�]�"�°���f���Õ��Ϗ��j�wP���e}㏞�P���l~���Ş�#NFM��|�zLٙ=p�Y!]��k'K���ɓ;�[��N�1{u��-������ez�ͷ���\�B�ڍw���P�>	:���n&�$�e���ЖRr�=�A� ]��?�8@+��nc�)E �{F�6�z�8�s��G7�jFt���6>�>�ؓL1Kϒ���:�aq$��������u4��e}3g����Hr�sk
H,mV��!�8)Z:���������,G�/�(Nޫ�44�3����A_�>X�o��}�����?��?{��Y��K�����Ԁ/>�rq2�@�X��s��L*�NK�)Ա{�h�^��1A�_�Aίu��+Eߝ��ɨ$�6��}��JJ�	C}�)�lS��NGEv�=٭������Ab�����H��������9Z�W���h�׮�w��S�ڟ ���RJ�5�/s��k���a�~�s�qYD@��E~���&�F���9�ۋ�-qZ��������//o4���<�ZtQ&'u�Äg{�!�lo��&X�)�LC��JR�t�;��Kn�˫���|7\�
.�`��KU����U�6
N��)���S�H<��49�*��e!�L0�_������z̾6|p�;�
S��=��I_�.���?~�]a4Nܸ(��Q�1zS=�WW���C'��"C�eS�c�F��x���m�Ff7�G�=ğ��4	�h��X��<w��w��E���kȋ���E�;��!�u�w�Q� `\�:چ뱇wo?���UY�P:�jZ`BY���O��qv�Ô�<z�#6�hY�
�ש�D�E�{�΅�0�'��ݴ�m���(��d�FT5r��+`ۿFTs�ΘY�w),r��N��tr�e`<v������@��gܯ��q�E[sJn�㈮��v���-�����=K�fcW�R��/8���^�����HE˳LLPӫ��T�F�)���
�i���%�ǈ�~J��s'�${��\�q��g�L��8�3oD��z�Z��:�Շ�o�T��"Ն�!��0�|`�x)KMIO�0��9���T1*�A?���6��hqH���s��۱�=2c��w^�t&6��⡥(�6=p����7,eufDuT5���!�F�(��������<�U�����v���&u�'���]�MC3���m��%u�-kNɌ�P���!(\=[ÅKa�����F�Y�Kg��k�J�	���.ƏE~�^�1��XS�}7�������Q6��v$Tݏ�M�#�R�����9"��G�=��3n3n����$Xd�j���j�P���/��m��Z�lы��Jǿ�|���Cg�l�z؎���?@�Է���m��y�v��\�G�[�G�}!Sz�BI�ЄL�7��#RVIԽ"�7�k�}�Y�E����f�/�?=�Շd�9��a�D�F�|T��������>��Ј�Y�5(�ittޫ�l4X���"������AO,�PVɥ��da�[^D�{,Ƣ���dW ��0��Qswxҧr3��@VYI(�gs�{T��6, ����X�ߐ��ho�	�/$���B�D�?�oįq,
k�Z�?��7��&z�E�1��۸x�*��3�wtG�����;�S�J������x�c�<[ҥ9�	�i#��<�ц�����`V�q�sU G��0�H��֖A����J�:��C�@�5����Y#Ӳ��Z,�p�-��I��;�"m���$v��2<d�7�/�>U��b{��]]ɱ������hլ�%o�����d�;��/1r���Cr��+.�Ʀ�E{��:� �9��Bw{���v��ЃR,��Z|M�6��WN��}������rk:}�z��ڼ��l����Y�������>���d��߳���5�Mj|!�@Q-P�ۡų;��5�<	-h�,K��yM8��0�@}͟� u>}�)�ME��`P���oz�-
k��:`(ix'F�߫�"""�jf��Ij"M2�B$��/��P��3�J]pC!�#���m!Mf��*g�?̍c1�\ c��!����xO�r3�.S�5��I���lRگS��.��N~F,�*��Sȷ�l�*�)��Y�l����	�L����{B��K�y��a[u=�f$�e�d�&FWt_�-�_|�X��8~Su)ㄎ�0l���B	g�����E�.\F����� C΅9������z�b�r-�RD��o��QDΥ�E��) 8E�b�J�&��69��T��~ź����KiCN��%c1G�<�F�$�ʬ_x��+v⣗\>B��z²ө�h|��� �,ƀW����3�%B/z~����]|i#U�1��)6B6`�}/�� 5����%�j�O�11$������yC����o�9�,֣Qo�hZ��@���N-�N�Jg��q� K
��:w��}b"\�9d�R錡�+߈>�R���kg��h@�|�$g�O��8M�K#J�V<��4�o'�#"�2���KFdٵ�S����L��/�ݦ>��������c�$`N��:���`�[lC�kY����Nظ�O�XMN�D��ҫn Ɣ\ܯs��A 3|]X�髎Y��,���K�&������Α9/}�'�ɭ��ʭ�Ԏ���N�`�����_�}��^/I���ƪKm�v�l�3�k�c�!�\��s�.��KЁI3�����A��2��5��vIy�Y�_�E̫�eIy?Ϥ�l�e�:�~`���b�v��Ȧ��ɵq�� �3�Uɭ�?(f��1�;���A�u�.�Mf�����Gr� s낙��smm�-t�Q����=e��S�%c�k�3���{.���������/{��=fLm��+�~1��9�2�Nc*�R�ţ��o�9� $�i,�#�rӢs����e�{��o�i��&}G�:�N;C�8�>8����G����d��c���ܿiM1-#�_I#L�&�UB��� lk���X�,t��d�D��lh	k���y]v�z�<}Ǭڛs�;CkY#\����}��gs�z=g��EM����V0�٥�Z�Kך�����.�g��x��c��^�w�q�[�*6�U]g�S�Ig���	Ȭ;C�D���?~���ml?T��9�gR���ǕX��-vQ��qU^"c4�}::��[��eɇ�D @�^���Xa�g~�
�g�����H�v�ݶ�N))���:?%��u��zdy��-QQ���`?ۻF�HC}R
=��]�����h��<*�D&wմ�U�Im�L��^'�Q!+�l���cQ���W��]�%1H�m�L�8�s�<�v��͜nk.�� ^ ��B+�-k~t*NWx�~����h��v�.�4�/a��9>UG+W��fz��F�#��˼�,�X�D��u>䜍$�o�up.��02ˠ��� ���4*�VW���k�*&M�;�_u�W��K�2j����Z�,�5Z�VKI��:��ԯ�rWCu]2h�pEs�xk�pW��4�-CyX��۴�r��`u����P�'4
Kj��I�b����`��ډ\-��U�YK+5�D�d�?'H�'�:8�.M3Jq�H���Zq�I�8�%�Ȕ��ؗ6�DӦ�W�k�Z��)c��g��Ք�$�\QΌQ|CN�cV��dZ�b�[|��sIJ;���W ���%J誌�3-��Z�Dz_3ZX�U���n4�B� ��U���`M3T�m���@��yǗ�ΰS�������¬�Ii g�30�@���9?���S�!�`}��\#J�Θ�l~U�B)A]/�3[�߿�j��bP�U0�z+���"Û��Us3��W����h9�+4�����)�*q��A�Pz�p�<p ��*$�r("������'�BѷO/�$(=����GA*�10`׸g��7�N7R���[N�V]�Z;�$277'�F	V)K&��<��_%b-���I��<�c�+qD)����~<�4h��Z/z'���/���'����C.���Q�yG�C�r��~��%)���ωP�%3i"P���!ӛ�d�����������#s�܁V�,
j��O�p��rԳ'{�q)<Ô{�rd-۾�(ֱ�y�i��H1�5
4�I�䎶X+�L*>�hue��i!^$�g���_nx�b��%:}�{��M���kO���h�0Pؘx��J4M�4���kO(n��y3�V>����=��L[]�v�j��z��H�U�Y&(�4_x��� �b�c�F�K��`Zb!�݉F&Й�l�e����|�a4��5��ajV�B�Ky]{�$ѹ����g[�Y�������x���Ӗ~�<�L��X���Zm��o�j-<��[�#;3,w�]���<�~: �v����!`,(e~�*p��R\�'��z3�>�RW7f�g+Qˋ��Q�<������6�fD�<���~\ś��%�T27�(���	.�T:A�ɞ�e*k*�Ů��Z3�TPZ����$�5�ݳ]l�gF���9~5=����V3	�ҝ�E�.� �tbR�xP�M�|��_����I��]J��r����A	�����J��Bt��^ނ��B�`j���dmm0}t��w����^A�_����q��~����sx�~w���2��q$�#�?;��� ���o�s�ƥ����H��[�/��Gp�U�x�)���H����r�>�S�4-��Nv���mE���-%�_#���5lX��~�{/������[������s�m��I��{��7�i��]�u� PK   � ~Xp>r�  �  /   images/c13bb491-011f-4ad1-adfa-58d33d2d83a5.png��PNG

   IHDR   d   1   ,�   	pHYs  .#  .#x�?v  �IDATx��|{�dWy��޾�~NO�L�L���<w�v���$#a�mDJC�P1��!N��ʉ���RvL���*Ɗ�`L��Y���Xi%����~?�{���}���힝׮fK�5)��ݾs�=���}�;�������O\��ͦ�o��&X�z]�д,��ʊ\|�WW�ihȍ���f?�y�Ѵ�a�t�6wձ��Ӥ7���}��5F��֩�ٕ�e�k5���0�4�U��|��;���|��ݨ5Lk�g�����\7�k�wBZ�K^����60eT�@���àۅ���fs{�R����é9�o���-�	o0�b>_ �j�, աNT�E�X�����V�����b�PD����h4갚M�<^�s[h^���c�~�jQ��՛�6���C�4Jyд�HLr��N�vw �÷���Z<_~���YM�K�	���)�v;͡��GWu��A�,��'hhfGnkT݁�_{���{�é�/D_�$6�f�r�X��O.\����+��!Ē��AAHoȏr�!T)��r:F�"�ȗ�Dm%Oɵ��W�3Ff����H�͢G~+�$n7<��=r��Yt%�omA����AdWV::������(
0�Qd����P�5��9?���1LNNbhh�TJ)caac��p�d�\>/�m����33�������A�]�ő��ҙg0v�8�����٩֞�d0 k`_c��X\ZB(�a�����ѣ8/s���*Bd��[����~�a�5�r��w-Lk�jqY���y8�=������}�r�C&�����I��N��jRM^״�M>�ԍg����(?X�	��X��	�¢�auy�,�а$u�#'�D�Úb���&t,כ�K]�\�f]�o���!%�7�-ܲd���O`�T=d*1�t8��A�yz�aS7Zo�{xO`I�wI����J���M �ǲ�w�u�	�(Ε�+�G0q��:a\�b��=�����cM~u�.�Wם�����(=-�(=,ck���H(�Ǣ�!����%Otw�+�S�)WED�X���E��R��S_�oL��	�h�Q#W����Hw�쒱���_"@�Zǲ�@Ƕ����Ւ�D:G��p,����#A@�4
Eda!��"��k��qJ̮򙴙�6��g!�+�:|��e�_�Z�)�隅��7��H�\�HG���.����~/���MIT�5�㽘ns�dG�"���
Uge�>�`9�����;�_NB("�]��$�/ͣ�;�� ��ea�Ӊn:`t��?�+�a#� �y��:���T������.�`w}8���� L]*��BT��^GY�n�(�J"�I&̺L�lH�ti�/�Pgy\�w�B�A/2�\���܆R��+��h*u�CC!>]*#�b]�u� �&J1�>+�?&<���%�9�]$�.D�C�n*=��Um¥GEĮ)��ǿ4Bd�Sɬ�X���"���ґRr� �VQ5Bm^4u�b�Ʌ<La�卢m�5�\zt%�A�[K)+����ҥ�B�k�糪, ݬ�QS�g䠔P5������S�H��Z�"�oʪ�69��]�r
�F`r�T�"\��#��(
���� 6"�ź��Y!�\���cT���-"*�O�HwXʐ�!T�9��B,�H6�b<7/�r���]��˹$���ɪ'�ůu�����k��R��w!�K�VW@b�ȑ7� 7ʈvxQ�6�zj�+��b�}[ܽ������BiM�%Y<�m	�P��v�ŏ{�eۨ�~�]�������7�C^�#�Mnl)b��.�����<r�q^>��f�,ȭ+1U��wMY#/�N�|.C"�%��-���K����1d������0ot��#9���=E4�\���LY��7�Z5[�SS�Bqz��l9P�Gm���s��(����^Dؔ.��P��G��"�2�gfWq~=�L���;-6�u�5ҏ�>��Q�k"��D�h"�SĒ��K��|#����dr��b�H4�%ѭ�K���(b"�'��-!N/�����|�{�_,X��"�\.;D��h��p�T�A���qE��tZ &|{�Ĵ�3�6����H�IM��fڢÒ�'E�5ſ��_��\��	c0��B��>(��/��U+-?����D��Y*"Iٖ�E��pA�����*Wip��Ҏ�2Y()C�����R9�m�p���"�0��*"+�J�J=����l�Cd����]���b�|QL@q�j&����+�p��f:���,E�,�b��17��/އ����΢�t(1�]�ؽK��hÃ��N�ΐP�[�5Zh$���j'կ�J�>���t�R�`�7�i�?ԫ�֒��h�i�z���l)u:}��ᑖ�k5��ۧ���C�ug��KMkY���Y�W�R�"?���U<1�Al�L�80s�
�h�Z"uGD��NQȤn�{�/��b�~"�H��|��e[�+���
�!ѣA�\���D��.ie]�¥P��8���Q�RH2���;i��)�V�{{n�������"\�.��B�N���C��bn-�����('b��|�4�+\�oD�}�!�~���2��v�R��!T�y��N_X���FS�Qr��2DDquC*�$����p�ًaKqP�P��2��UAC�ԪR��Q��]>����Fw+e���0�CN�3���];�p�Dφ\���؀\�����0K���$�?��$R�m���Y��h����ex�������w�Ƹ�>���Fb��E&�.0`}�Q���{����������|E(�D�X�Xҡ��Ԅr���sgyI�w�E��gr���ƺnᶁN���1�:�8���Ȥ���8���yg5W@SD�߸Z�փ�P&�Y����$��iM��'�)�ծ�!C������m��CMGQ����:)�˵ֺ{�%�-��s���xj&g;}�(D-���'���.�wee�1��ư�ɪP��Ӌ�5	�Y�B'�P�ni�T���4�e���q̊����&>���_�G��uEB��o�#:V���cZ�coC9�#�!�,��3�Ю�ZADR4��ٲ=W��i���7{GGF�$�/-��4�J��L�yPG�笋�,�v!��!��V j\�p�GS�9:tY�+*��̨�-�t|��wQ�����ĕ"1�:��)
�n/����0��_����=Jw��k�wcp�%
ZEz9W"�q�h0���~�ד8���tFE�a��b����8[�G^(9��{h���ͤe��H��Nn�"f��fE������;fz��=A��r����ZΥ��ٻ]d\W�o!��@"1��X{��Xz���_?�B�TU���ۏ���B�CH	
c���jc�����s&�EMĘ������;;x���um���\Q&j�x�j]��5Ok��ɺ�P������T���&y���{@D�p�6�vw�60��Gw�妎'��P�+xO����ps�I�D�q!���@�܏�?}�P����ٛ�c�&U�ײ-0!�r͂��|fWLr��"i�Kٱ�.J�p����c�i-5���%�uu$�5T�oˠ��H����Z���y�a����
��K���r"��f/��	ȶ"����_�"����R��-T�4������J����/a��3�'��s�����sO鲥�����Ṅ��=�n^e����B"H�D�AK�&z���^UO����"?=�Ӊ��2J�+h��=�D$��H�����u��{�@7ַ�j��g!%o�3�j�f+(�"0];2-�.����8�_��_�ן@����)��!���٭�%�^�ήؖ��3�!�b
c	?�s艉�0��3��(�D=N:j8�яb����cڏ�~*��'��t ��`��h�o�nLtca3�D��,B����I6`uD�ٰPsy�����Eyg�TCI��)qdoL����&F�!��+�w��l��ld���GQU��~�u�\8�l�w�s�i�t�|f5�G^\���k�����3p�8�?�t�h���V��� ���T9
�$d�+G=dk;y���k��فB��V�3j���johT�-k�R�P۸V˄"u��K���?8��ׯ��V�t�զ=�J�ڈ�\N1{˰�G{�Ss+����x%@�{ؘ��RP5���QR��f�f�g5�E�x�62�\ �r��������N!�3R*�j{�~%V�U�zl���w�������%��'��3��Af�t6�̨|�JD�K�q�C���yԅ�F�r=�v��2_�b��k�xS�0HX��Ⰵ����c����RNcL���x�ٗ񫷾�x��s�G����-�".�9��A����<4ػ�*����"\���Ԣ�lq׸l7�ہ�߇�D{=���C��^�TɁ�BH]fq{��w��W�XJ:���k%����5뚋-4�8L!�:�~�����x�,��I�����p|H���_�����b���݉}�[
O�.�t�T�,��WIps�J�!��x=�B�ob[��j���1����&��f/�-�Ft3&�!�nx�`�fY&4��u���ģ,�9~J=�v�f��'^��>p7�ϹY|�k����|����8��;nƽ_~�r�8�K����p�/�ŲP/s�j"��N��%#\��D����xV�8n10�]�!�{�px�������e�n��-��>��m;D�̕-��ב�_{��B�ܩ��_��������o��ď��z�Gg��g2C�p#�]z�B��i�NzA�S��R��D���r��$U�v@���]Iؼ]�W/V��;�콰��b�rx!�_͛��fْ	'���,�������?����?~��ދ�gV�Ȣ���K_���v<��ϫ���~�x�sxaa����#	�[M�	̹�Wn4�)����Na9�)�[-�R�PW��S�s����ѦL�V)R�Y���Ĳ�ƀ��;l��j>4s�̟na���ȓ/�)A���.��K�
1g���R��G;����_S��4-.&Q��>h�������ž��>��*�O")������Q4}����%WV+��6BFGG���>���U�R�v�p�L�z���Tc� �ɪ�+��`23�#`|���M�w�x<�+�P�=�kT�T��)S=��F�SO�,H8=��R|�@���Q���9(�n�޹E��xw�2}��B��c���B��$�����zJ�8Pdu���`%w�Z�1����@�eǌ��ۨ4�D�k�����wu�pa
���na��
�=:N����yL�����{'�VR!)��N`�[@��%=�ɍ���=�Y��'�vּ$�䍩�dm{ϝ
����P����f�w��XIe��q1�W:y��G�����6��M��tv]v��Xˉ�<��J,ߘ���>��8.>
�|��_=�WX�D��~'�ٯ~�H�|���xdjf��>Ni��:LQ^w[�Xv۽�gD�������'�l �^�}��JK��6s�9ж׏�8���,E{�5r'���~���uյ&�guwv�:�p\\<��c�j`u�E<�O��N���6�ʶL�����-<����S}�puA�?�'����W�X�=DH۟Tl�j�۩ ��]��@�L�ǽ�\�������m��I}�q�cv�U��C�N2{P��$N�N����;�<U��4p����[7���(�Q]C����alb�Z}�}l�F���au@��	�D���S�[h�Evg��X�k;^�^h���V���g�-��l�5���<o��3�e�>b�,vZE������C��+����7���9s�i봕�%
��B8UG".��P���JU��fg͖x!P��*Ң���ZU��#��"��Ib�����e�E�im ���X�u�p9�9z��c"��
��ф�:cC�D�`GH�!x��f$��iJ�ch��b��m)hM��Ʒ~�[>4+>�3s+eC���}j�-��$��u����Xm���1������ut��^�BY����7~7�����{���+����9@��9Ãe#�O��?��֖pPC(Ɖ�x^Cѷ�7�;�%\��i�l��:�H�sH���::@��0�G���Pg1��b���BŚB<�M ���c����`��˧_PQ\"�ͥ�9����_�
8�o�)�k��?�Q?��3�U�\2�4�,�x�u�����s�>t�B�erPv"���:yD��{Q��DlY.��ݨ4�0B�B��ya��0�=xy�������BIwb��B.G��h�x�R���G�\Q�W���nLt�{���Xr���S���ʨ��J�0��y�I)~��� 
b��Eɦq�/���g�j��2���Y�C����s�!ļ��,ƺT�J8�}.r�UǓR.r.$"k��;X�xW3�
w?�<��������8�=��Zωǿ!��K���Mv����� kn�d���g��Z&L�����$4� �?�a�6�ؠ��,S#/�V��z����Xb���i��>��#X�[E�j���E���\�����1��Ry��|��re|~�k���L=�`�k� �{Q�)v�2�a�X8�tY�/���@P�s��5�)8�K.>��yq���fϟ���)�(�|���3�#��x��C~+� *�]9{�,z{{7�B�V0,z��#��5ܘD����׿��:1�(�n�XvY�-eZ65���7E��=�Μ�	⚁�|C>~���~Y���$�g�U�~lȽ?:�B0o9׫g�&�v�n� �����
�צ4$H��v_�i��H0�؄Lq}�!Y{�F����9�N7e:V�ί;�wM��*�y}2Nv����d�E�땺��R�����`#z?����
�-?=��d�x�r�umy�_]} ��'7;�����o�F�[��Kr������l#�`0�B����pH9K5��z��133���qL�o\X��)�1��߯"	bũo����9gRI�~��ȅ{୉�|����p��������a�$򻾾����H���e�����o���j��K����4"wߏtt .���a��2����oJ�7�g~[���)�_G�Mw!;J�~E���Z��wO��$a�O�8�t�9r2�jY���K�o�5"ױ7~�N(��1w��v��0��h\��@�1��C �DL�����[�E��:�N�(u=�a1��� ���f�e����(�&n��*��qՎ���G�J����N4�.�W&2���8Rސꓙ�������/q����R/sxk'J�n�$�1Gd������/ɵ.�{��F1���*�\��%�����u�\"����lQG��	�:�0�ힵ���j����rw����i���s��#�8��wn�~�Ĵv��m�s�:M��םb���M�o�8J����n�p�Q���:j�i�*�    IEND�B`�PK   � ~X�+�s;  z;  /   images/f3037bb0-f56a-43e4-a2ff-17056f7c669b.pngz;�ĉPNG

   IHDR   d   d   p�T   	pHYs  �  ��iTS   tEXtSoftware www.inkscape.org��<  ;IDATx��}�dU����z�B��=��ff��a� E��~���bXu]W�[]W�.:,b �H�!ϐ����=�=�su����ι�UuU�V�ou�Ztͭ���{���p�S^i���6���-��d~���q����n�%�c)E�Q��m2i�΅��Xi2S,��'m��.�FQ���-���Tm�����b0s�;B�~����e�>'Ax���;hW��������߾Om�P�-����sC�z�C�"�"�ZȐ4]PR
��m����5�������(|��D�>u�
e�ڶi2O]�m��$��0���9@m�������+��XҰд�OP�1,�|��� ��r�:�P�����:駙9E�)�3��5Pn�H��~{����mַ_��|���O[�)�٩����~qme����
`q���eIm�ō��!-o��/@Zє��7�dڶ}�|���m�
��-��!��he��x��u��6�o��~������_�$�.Z|��/LW����yf�!������o���h}/�|s�o5$��`qQ�)^�Z�,�̲��n�V4��8Ǧ=�`���e��J4#f4���`ZNѵ�iM4�h�Ry@��Y��3XL��Ч-F�����k6���,��LW���a:U��!�����
�<�.�0�x��N詔<�Q.�f�dw@���H�t5�C?z�v�f�ॕ�g(x����sYRa��]�^��Π�)�Ѡ�fF�Y�o0��C0��+p!�h�Iv;�H�8]���՗
 ڟ��h�4#��H���A<v����A2ɫe�{��caV(�(�Qiy����X����3�W3��@X��?�EI4c��j!]�"�� ,d}�D׮[涯�xSԥ
�3�2�b.CZrbe,�2i#;}Ƞ6�d5k��x�X�F�`��h�o\i:㼹�o�K/<��4�Mc6�*�Y1�g�b�)�L��E��>y�يܺ�652�=/�P�mWHa���H� M��Z
3�3B�����h'K*Mk1\��cC(?z of���.j�X�d�X/�Y�Ҽ���n��iE���1kD�͊��u'�_Q���n8��c�n0e��ym�à]2��ߊ�T�u��=��,�~O;�;=�K�n�"V�G�VB�zR��GV��D�q�[�Y��[.-n���Y� M���1�%B��Y�R3���������Ĳ&X)��X�X)\N���8��������{~���*��X��4#��j藃B�dY֓�P�6�t�H�����f�̥��>�Į�M<�U?!���|�}˜϶ؙ��<�����6��p҂���nz(CT��>���]���߲����[�D�چD".�a�.�߇v3"�8!iU��[ݼ��4j�9����#�x귏����c�觕o,}~�1��WRʂ܈�4�m���$/Ȑ1�6�������ӏ?��J1ޱ��,�u"1":���L��qO�Ik�Ѯ�!:�PuY1��+#1T66b� �x��)�E�z��P���ebJ�p!�BMQY5�=�@_��y����s1��҃ŭ��՚-�]��}��`�Lc�4�E1�8�hV҇6{F�+aAMezN��J�Lo�$�]]���u%P3,�)�c�D&����&�������D��ٝV�J���54���[`�B��2f�V;m-k5�uz0�?.�d��8M3ᯮ��ӅvR��OΨ�l^����C�3���'�(�Hf��,�o�&�^�n�^y�;_�n5m��F<���*�d�[�8��z`��J�`_��D��;��!��VRן,s���@g��p8PQQ!��O��eg�����)Y(��;��o�.X����ΚfX��0x	����k]#�k!;w#�3�:넥PK�C�`���:�E���=S\\�?���H*�Z���Ls�K&��H�h%h]ؾ�!<���(00�L*-�|1q50	}�82� ���X�N����o~�
�;C��W��";f�A�Ě�O���P�a�>2u�R*QP�c+t{0��|r(�F����f�ʈ�g6�^3܇�ۿV[�\d)n���e������Շ�o�C~4�r��U$���i�%I�T���좉�!��:aŮ#�#��Q�%e�����E���}Q�����<�h����4GؿEE"qv�ˎ3��B �%s�%�/- �3s��lᕖ`+�f=+��i�\f����P�I�ξ6}��-v~:����-�CH�&�|���{&Q�b%�z{�EgY�:����:������m�ɫ:��x�x�w�'���]�ǡ�*�t|�܍k�����F�UR`��K<��[0����o��zW�>QgGR�����'ahC�=�ъZ����Qd"���z��ƞy	�?7	�Q2��C&6������ߠ��sz�p����.���HX�2q~>����Iv�2ы�Ƣ/�'��g��iH�;}U�V�
��t�H��)�����0r3C�0������$��̶<p)�m�o�9hi�HN0>{Y�����E��CB�i|��jH6R}'�����4A�kj�*L���V^)�(��a���O��@�k٢�$��5@'"9������D°R{=Grt �8�d��Zh�{��TYEmbЏ����*�4�3�K�ӥzV�Ok_h�� �B�A�C�n��g�gƆ�coB��Y�����j�7�L�����	�W�L�c�]O���m�.[����u��P򳏣���a)��؝�G���!����|U�y��ct��H�1$b���gP���g2��?���J�$������-����v���'�p=���^��@/��%p�{���;܏�+އT�a��䋯��Ӆ���,�u�QMe]���G����:
^�!=Ǡ���#���,�C�����X�H�UP�e�p����lM`5w�.\.�f
7N:;(�*e�I��I#�JqzR�}�t��S��B�ij�V�DM�O�����]�@�O�~S�Q�-�
_K�*�O��Y/�Eu�?�pԏ�6�c1�%��t�sa<�l)�bvH�woC�?��.+��4�.�i�ҎE�J�5��@Z���"�=��Ϡ�̷kl4�IHU.���v��t�LP^�R� �i�T����5H�hB�:!���	!XH�����-��ό�BO&��0��#6��C���T����a�R����Ӣ��	Ȓ�>Mb��!{�P��nc�)�,>3$2��i�fxኘ�0(Ғ:Ns;q��C!��yU���S�c�7����k"@3 ��4�ii3S�y�Nz�J�X��e	v�"`�;���:�B��
A0-A��;��7"��FJ��H�B%]1y�� ��Ĩ(\OO�c�G���DL��J�[�x&�M0I�F�X�'��oC���n�`�D��L���H��hZ��	�}$@D�т�1��y����|4J$#~��I%��f�"ZS��� >�>��UM����f����v�_Nm��5<��`�D�'�UX���H��~*�#�l��*����C�o<uJ!fRC��0�K�����Y���ob�F����cV��?�=�x��&��e�~��%=
3#��U^�:���ue�8�)"��9�"��b\�~9��������i����7�?D�_nw��M�L/��M��s���s��9;d�P�=�O8V-2Z�du/FN ��_/�ȱ!�0՞v��}���%Bm��ϬϨ�0�zF�N��GF7��r�i[8](�X��uE�������$�����O~�n9c7]������Ӷ#��au�浈%�L�o�Z�E�$&�7�N�Y][��HN[��� 95�W_��	��c,>�N��w�����n�yYhln�燈����k���Mm��a�/&�Y�q=�B�lFt��z�G���0�g��9�^���f��� �iaC����!۬8���9h��=p8��$@�
��h��K������o����VU��uo�R��[i)DШ��d"���
�k4{�f����@����Ց4	�z��ڲ�O�'�E@����MŨM�\�v���k�ꢬ��xt0���T�(!�p�ظ}��CH�;�g�����,����K���Yh���!�ӱ��t� �L"M%�CX�*o>�?��C�y�dt6�����ק����g����eE�>-���/������x�p$f�8����ԑ� ���Ț�!�+��	��ʜv�=Dv����N�|�KA���7�B�1)�ljNQ}�=��;d�!�H���3��=���@s$�K�feD�f�C$FL/ll��;����V�<��7#�XN2�˕v2jB�˝�@�����D��k:��߷dt=Nl�p��\�5&�tQ%{|S��3C�sP� Ms�Éd<1�������d,mY��7�wS�_�wi�w�4��~�~0������Oi�Y4L���%�00HD�&R�F;�s�"����*��;�}���e����v���'F����f�&�_}��}�:�Ēp��������n�IcwN���:�r2����l=��X�픭��２�����׊>؅�������쇢1d����1r�LzA#���(�"�P�u�[�!,���сa������rܰe�	?��r�B;�Ey��a9�t�cU�;ػހ�؎��!A#�$��meY��s�5@����2$�	bH�]2�t�1c����\=�	v�����;��=32$�}n��a��ײ��}q�"��8��
�{��@������1V��@�4'8Dk���o���",;��-ȹz�����:�A~��ާ龳�!|����v�a�/ːI٭�myF�$��bV����b��w����A1CF3Sǿ����
s�'��?%|O�Oe*?v��fq��e3����-4���F{���>���^�f�_�������2�nN&S��=��b�,1�E�����F�B��b��n�Ӥ/��a���r�v�z&^Vp2\�2�'Ơ%�0Ek���ԊL$�����Y��U�����@g�^���#�u��{��뀕���2�#ƭ,J�}Ub�����R�B�׳�a��HRȯ��"���J���$�����
C_�sti��2-9$�)��UX��k��D��vH�D�}��C�"r
e�\���F�H�����.F���_q5��
��m@��qq��K�@���&�x2g��E��h�_��I�\04W)�Vݢ��(�{(�� �~qY��y�~�5(�{ 0=��`��P���pd4��ë��ِrb�x�LJ��W�vHn��gZ���Đ�e5,En��ȁ��\�$¿���h�I�7�#nm?�e�����]t����!�~z?�'3��hVL��(+�'�'�![&�Q�����PgL�f��~��AKP�@.f�Ёي6[��\�~Y��� ��K��ٞ"�'q�z����Bv:Qt�F���?���W��l%2�\3�r*��������)l�횋��&
�b�|6��٢������I�e2��8�W�2)5�XA.dk�������0���,>�\�[�b�W�@:�l�Ӫ�8�!C�.��]P|%P#!�D0�³(�~�����
{0�QKƌQҴI_�@xYhN4�0��� �(%�BɆ�z��"Y��j\ͫ���#��+p4��:�t��u#?���V��?�A��v��(m���b���#(��5��p��'VW��?$¶��8����Dp��g!�櫰U׊	ȓ�VY%Dw��A�ܙ0� ����m�VQE�"7��ar��L�@WS�@FB�Zb$$Y�s��1A�Ǎ�l�8w޿�E37N�1	 �z�D���C��XfxXYXD�XQ��fأ��Ӌ������G&M���`	b�ٽ��	�[��i'��:Խ�dB�GM��ޤ6g	z�{�i��썶��iO�<t@(��Ѐ�<�N#������V�
���;���$���[X:�z�ɈP��(�w͜La1�Ngo#�#@���pVz�a�Y��ٵ���2�cN�هk7��F��wb����U����H��B+�1�� �1%�oG���D�o�V��.�/��s�a�0_�
�e���3�Z����d��ayE3"yi�y�V��AݎǬn4�^��[����E�"�cq?~/��2:;;c�_V���w�Ia��~<m��Q|݇�#�X>�vZ��|�k_�/cC��=�1�G�B7�T,��A��r(ⓗ�gl�ǯ�n�:&,Di#��L�W�G�n���?�{�)���"Z �a�i��amA����Ah4I���'�4��p䅃�R�(�P,L�J�*�|�g�A<V�̄��-�i),�憢-`e��f������^�+.�^"\6��g������><�������L�1�q��V=����i��W�{��N�����&Y]L���$2v��D�B����C��'�Z�] ��
;Rezv�W��-H?|nR��6!nu�%{�T8��=�뗠{Z!�H@=F��ƿ��+�<�V5��	�3*I�S<�[u��ۧ݊+;����DҒ�2�� �ǘ�@~G1�~��P�?���9Kt8S1�w���x�[��~��⋌|�drF[�ۍ�r����b�)fw	�X�f�Kb,��C���aܶE��c/l�r��c>�b����!��C�¦�{�|��HZ�yb��V��p�57N#}L+��9,��}R'��>$��ܷ�����k�M������ʍh��M��'0�ė���-���3O}�8�u�pa8�"1�����%m�`.�p=3���'oڄ"~�9h�h�ӆ�n���>M�L�q�	����$��_R!]��5lw([�>4��<#'�K���6v�JvY�hʆ��
��꩘^6��>J����U��'�)�$%Oޓ"�y�Wx`�bC�V��eZ9�2��-�W^u��\�(Y@��сM��b�E��х�9�f��!M�C����ڇ����a�V�qZ���c�A8�[HIy��@�	B�_�S^J�,C3K�Y�E+��bS eǓm/f�*$�����6��d;_l�r] y!��?!�0����g�M��9�4pk;w ��DG�+~���tE#}�o��+j��	�� �(p�%^C�=.�Sߘ<�@�Y7Ŕߡh�W�ؐ���%
B_��͹�"[�Ղ��}E4�{C|���p�Q�dВ1X\ޜ��=�(j�:�&�XYY)`��~���	/��"�2CfIr���`E� ���F��w���;9����p(�7P7N��,%���ɺ��pVT�}�K-�U�\�>��Ŝ���0;6	�{��%dx}��_b�m/�ɑc�����,8�>I�e���R#1����*w�\(++CMu�	j��̙���ƻW�p�d�$�h�����'�R(�x�ڍ� a�A�rF����ņ���`�ß�{��<�JL�~�= _x"0�
N"�ԣ�#_DQ8���/��D�\9�+#!�]�E�2��.��d���
��p8��H���c�/ Or�I[,EQ���x�C�#�#�%��=�Xk��bt�0c������5t�n�v䈱`��K0U��g&̸'��tc�3��D��|����(��:Ay$�e��хzlJ+�EO���a�H�����pCQ,S[60�i@D�0Y�G��!f��8󯺺5U����#����h����Ç�q��֬�v1��*2��xb���21&���o3�~�, ���֞��}�8�2+�زb/J<L�4<<Hv��N��*n�?X��"�,p��!UUU���LQ$=I�B]�BkɴL�k�	��-R'(��D"�λ�����+�PRչ���l�%.�,���B3���hoG�"C�|[+�o-��V�sX���&e0���{:�%��԰̜?3z�V�ɑQ\�e+"�Q2��ˮ�h_m�ˠ0[U#G��{��̲"]ŵ��7^Ƿ�������[��pS�EL���FaUk�1����ۈ��|I@� [�Ծ��ń�M���[n)@YYg�0������,1��Ċ�8ғC`��۲
�S����E:�B�Dn'��GM3�FY4.�ˍ�d���Uը��Ĭ8���	�&�U���f��b�J7?���d�󷏡`7\֮]+c�I����}xf�s(&��,�l��l�㍞�4�5��e���@g�S"��}Y�#X��0���(��*����`���;	�T��d.I��4��@� ��P��]������8����F�57>�������>E�8�����Lx���!�Z�
M�a=�H�����µRc�#u�PS4�Uh�i-z������/��T���F��~�`��b�ϋ4d`` c��|�=Z׬1|\s0�Y�q�Dx�wX-� A���7�N�I���	T�!�h&O�m��+�*��[s)uj;��Иe�p�Y%%�������8�����~�H@�0S��q>��=�^{F��`k��\B bU�z�n����@U]����
l�Q�����"�W*.���D�*u����&h��D�z���3W��4F:�	x�⢘|ԟe�n����*�X%iى�{�xz8G�*HӺ��j�n���2�/L�"�Yb���8�&�M/̈��^�S�I[�I���ҁ�"SXI��e�S3F:�}�#���	|M9M�O{��]��4S�؞K�еե��|~���9��4�	�zpa�	����:��'�Q�NzM���l������.f�[IR�$�.�����!�zc^��Z�
Ȭ��ŃH��%f�[Ҁ6��Z"^��Ļ�}�S�np�EƲL7��PL6�H&�Ԝn�̭��s��%9����"�W"�����>�n�B�m�&l�&��<Y%�c��/��ƅ$}�<76���ǡ�3��7�� �Ua�I�����~�N6��[�R��a�<�^	��):�O��}8j+B�KAM���(F�:�*m9^�n'n�����p�ھ����Ӄ&E���2�W#zp�'���ߋ��h��ۍ`�	|��# ?��ag�x��Fr'!\'G�n>�p�x��L�-
��FFFP�~-���j�oWz!�IhW0~��aTUV���6��MU��?���M�Aó����7X�В��t�3���>�I��`�-��a��j���c�h.;����a�:Y��e�Wxx?�������=d�0�a8���|�)A�އ{t'A͙��YtG��Q�i"
;;N��|@A�P&��:E�IG�<St�2��|4>��b:A�k@(�0��DC��**��r/!}�z��ć�,Q����O�O���&K}�=��1?�)��p�s������y�#�8A+㹗;e�w;Ĕ���G04�4 Y͹]�*xq��Z��>.ғ\�Z=|P�K�rx9��l�_ºj%��<���ݹ�!|E�D���"��Jp�����&{g��{��9��� w[{��}��dk:�O�'��
�A���A�P19�uB��đ+pP��JJJP[[+���ȉ�jG�E6�<��|���R���&�1*�d����OJ�.H�z�
]$�͟��̨&��!�:Ja8hL~�����;}�L~?�L��3�!��8qa�'w�Y6��#�����_Ax�F��4�������L4�e�턪&V��k��N����Alڸ�_v�ܱ�>�(���66`���@��.�9b�X}%�^?��W�QRQm�(
�$<�.!㩟�ub�h*���j�e���+���#�����\e�����E"�|�>LsJ�M�c/��.,��`I���C�xP�_�au"�X<dHB3�Kl#�"�;���՝��34�Pz9M�Ёɭ�D��Kn�-[�o����.l�$�b����[�ك�^Z���G��P�����=�z��`��M��T�JZ����N$o5:6�[O���}b_���+Ѵ��h�x�U�2����=e;��,�d�`Ög���[C��~�$I݆h �FZ�	}3y�\YfH�~��L��$N�<�#�w=�����Σ����w�p�͂<�椩�oooǦ�N��%�}��b�5]�ޯ�iSv�p=�ů�g�^{�G��}�qU�r,�4�e�d6C��T��6�uB������'D���&�E6���14�M�P�#�1��*���g����fiqĐ�-�səL�����	#���iF�S6�['tF2�p9{���c�Qݼr�V���C���x&����g�_��ݮ���\�"T3��=b�o�8˫q4���چP,�DA�a�l4�W+	\alR��#d9��������:>t@���"�Y٧zc7���jY���Qw�����8����w
Ĕ�;Q���Rz�%����V��N�(Ny��{�J�uv��!v�gl�"�w2��+?���"�/kF�nZF��>�Bg��\�ؽ�m'��ϻ�x�`�F����� j�����
�9=ة{jjs��J7-�GFe@1^8A-i�1x_��&�1-��3�5�l=KlSQL>�4<��F�����M$F,(jY�T_����G2)n�8�H��@O���#�ۀ�@|g���+ϋ�
����!nK�Y&E޸|�����>�gt����Ҟ�獻�%��J��)���g���:Z��Hϓ�i#��X��o�.i�Wu<��,������蓄�톯_2��L���[$sv�M:jz*0�\�;׵""�<>��\,E�[o�,� C=��C����aD��`�!��@"��BǏ�H�y"P7���u?�G��pM ��S�˼�e���Fq�v.Ab�cɮ.���n#��!+���6\�!�^���$&�T1ƤQ�;t�C��=C4=��+���QxRQaq�R�s���=�:'iZ���[�l�d섽�A������u(�����dMK��J2�q�1b^�9����Ȟ�#�W����Қ�:q�
�q��%��O$MM�ά��i���x� ���	z�]n��WP�U���v$����b��P �w���%w<�˗§�IZ(�+T.ݶ��v}��O��b��^MR"J�]�+क�	؊��4{ݰON�E2:v�؎�&��(�B�f�N�׹�T�[OB���H���-kB�d��\�lTo1ĥ��2MԨ��1�Mے͓���0c�o~9p� .��,�P�n$��;O822��=>�.���J�:W�3!r`/�$�#���ZS�T$*�a:[�����!��4�Oı1��/�U�\���~��.x��Ι����v�vثV������?*�Qݼ =|5�����q�kP^���ŞF5F�՗s�#���{ϫ�QG��b�J�J��-^�3���J������*D{���E��R\����)	fV<����N������b�����"$߽[����w�}~�[σ�3���?������>�?R҄�n����)���	f����[�
S,���'1�%��r��r��mr�K<��r�6�S�y���c� 4;$�8X�<��� 0&i���?Ɨ��c��|���ouu��F�ܫp��X�Q���h"�,��+���z߻Cl�)�~´J�6��!!N����9
�(Ь����8c����/�燂�V��Õ��V�E�
����bqó�\A\�j���&�����w�,2��kk���l����ϣ%�%`�d��0�����!>�����y��D'�����w���s��>���p:��M����[��Zojj��3�YGɱ�����[k)�+�ov����Q>6������4����غ��<��X���-JHS'�H����Ŝ5<uޡ.�ϲ`�D;���`ǵ�@��Ni������POn�c~"C�H�ߣ-�{xX�>��?���ċ�}%#����
��8V�g�Y��8�ÿƱ�n|���ओNY�<Ax�d0�ǟ~/��Cv�W�ܣ͒�Ęs��/}5�ӳ;�����5��[��}��nNv��F'o��ྀ̽s�y���H�Q�;=����[}����H)(���o5�!��J��H�1�ɨ�Bh���0"�Bm_%��co�����W�2
�3�g����뱬��'wubt2A"vj�q���"S�"�p������GCC�4�]�������H�h�T%��&5Ǵ�[�DL�N�\V��V��kO�ˌC�/��T��N�J.��.��|1���nCI篰�p�8�)CW���KkE�n!���`�-��Ѩ084�~���wC�"]B�L���g�j��z�2�#�ܗ)ű�w@"�u*�0���7� ����2�f��ĔS��X�j� ��{L��s-湓�D4��]9�jxz�{F0H�т$=��컛&�
p{��Đ�׈�-�rbf�<x�o�ג�'S�֪
�%xxx�ؕ~୅�>H@`�.>���"�S���Hv���a��˅b�/3؉u��u�p�}⁹�����ԥ��V��Hb�}�rk������$#AB���1O5�����n!)Kbq��xN^�Yc0_�����Z*�X���l�t��!��.���^ ����rb�˛��ݐV4s���,^���&^��o=.H�{HR�y�Z��� ���9�u�J7�у��Z�hʐ��م�"ZeV���4�d`n�Ԍ5��3b�F��S��S�� ��E*?G���P������˦��=4�Q�ԧ�:D�w������01/.[�=0:�	������II�e����i!>�ה���5��$�1E3�2��դ�V\',vf}=��+�C]���!5��!J��o����^%^��o�.|}7�)%�'�@�h:�}�=��P�~9;��_A��ԋ[x�X"�X�J�����I!9����O[����@H��,����Ѹ�L$11a����,����pd҄G��IBN���"@F*G�,�XWg�{(,��܌6�y�t���Z-	�$�+��_�u]����Q��J�af�n�b�rb����Kj���̯�f��9V�"� ����@?�À֚��Nf$�)��03Z�u���{8���&ie�=D��_��H�S��Ey�6fF���A��/6�#qw�/g������z���p�l�ĺ�:���rPkYC�@asÝ�Ƥd�hξ`�7CK���O����<j�A2��Vd72�x�&o���k˪�%h�U�S���4.�[`#��&�z��T���*¦�H�z��[@c�j<.�pXr�}�b,	��������mB)zV��.�D��{Ǆ(.�C%=8��Wn9y-�����`Z�����eZ���gosh��R�MZ��!ۀ7�Z��;�$⪞J䗳kO�f����]QPJ��C𰴴T���WI��'�$���Cq+�	11øp�>��9�<���J�-ƓP]�VA�ׂ��W�U�}N�Q'�l�h�NXeS.��"��yC�@Y�?ہq\��f?�z������ET1�.o;k1Ђ�>CY5Ը�W�;V�-�O�<F�W�31�ҿh�2����}�����w��V��Ob��^�$��I7�����Dk��ܲn��د�DVn��n���K8W�&���w�Wހ�<⽯55�Ѽn\�R�߭��O+���B(k��k���r�D�-����)B5Y���G�[i���z�O߄3�p1ڡ����E�YMm%�VTQ8b����X�B*�� ;����I����,�Be^�'z�i����l����al�#��<�.흃�b����q����
�r(�t2t�3���Ca%[G�ض}ݍ��
.!yG�u=#�]����~X)��l��.o�U׊�B�3��S�.e�H�Npr��A��$�O�/Oo�K���P���	G���=�����xd2��[��U)A����C�2��e\���À3������$z��X�:q��d�P^b��t� ��G�f���V"�d��#�ә�+ԔP�)o����K���7�k�"�A��~�zACS���$ho�3�q���.~��KjX~/M��km�E�pޣwuؤ��c�W�V\0u��� ��IؿV>��V��SCp�+��2ـ�᰺G���BmGt�V���ŧ�,��&nk/rQۍh?8�J��S8�����ʋ�9m�� ���D�~"�l��E�E,�~R�c�e�H�ץ�Շ,�ʺ<4B�.#��M��&ɻI�3����Z���v�b�b�c$	4e�eR���5��}�m���~6Ĕ���^�i_���O��Ж��fb�&7y����c�g��$z�Ľ�ޏz��`����#�ȐcCLl�5N���ࣻ����bbV1��Lz��ڲ@R��3�1s[��m9�C�k+e?Sǜۈp�OL"�A"vS��2u�ܘ�D:� ���|.$��䤱?�&�B�L��mMNX/6��2F��ߊ����@5ι/���Ǡ�qz�S`9S�C D;FS���z��&fӜi?��|�-��?�
��m.BUg�h��AB�˃=�q�]x�tG��T�����q�\�I���e��c�i�xz�lgP��|���ݫ������� ��D��s�F��>z�7��Czl����`�&N8�','g�6�"�2��wb��;�hX.z��2V�|H��������>�H�A�h��]$����cF!CL�0��G��,Ѝ��^`�Wel�w?�'N�	[f�s�0C�$�rK�� D@�|Z�i7�9��8�ϫH)�%��a����A"f���B�4r��"��Ldm�=��OT�zf�qĬ,c���}�"�ħ��~3�x�
A�,����Z�U9���.��b?��SH�E<�h���"\��8�%���.�i$#p�*�"��
�E�!�sz�ԣ��	�=���d1QO�W��#�uςl�S�=��Y<�.D2���ȰnO{a�t͖���o�-\b�    IEND�B`�PK   � ~Xϵ��@  �2     jsons/user_defined.json�[��JǿJ��]m���2o9���#f@���V�m��R�NB��~�N8�%@��<�����UWuWχ�����/�����]�v��/�oݰm���\��v_��n�����͵���}���+��Ψ��_^ٝ{��������vC�^�a�r1�[�]4v�u�y�_�7�dT"�CFP���ZT���/�}��m����C}��y[��Z�-�p
#��E%���f��kU���]�	�p'��pq����i�ˮ�����~�n7k��q��1�����o�w��~x��}׾��!u�����z{~V��m;���]�OxA��E�]v��~�?�_솽���-�x�峛'��?.�TRy�z�r��X��<y��6�e!V���%�<�*T�%�"dj�׫$T�P��P@)A�.��PB)��I�	�����I������I��PS��t��PQ�K���z���_�44����R����(,��*����PP�&Š��V	%ŀ�OҚ���0�IZT4�?I����b@���h(+T I늆��f���%�^<~�F��\B�G/V�4:�1D����L�E�Ơh��6���B�j���W~�`��@�r��f�,�@�?�`X$�(��QgБ��h<��=��c�4U���ȑ\���49��ayr�H
�ϓ#�$T5"O��P��<9RVB���dY�i#�<9�hS@�ɓ#�6	$�GG�n�&ytdǡ�yd!Ǡ�yd9Ga��z��"$�]�V�<� �0n�>����)hD$�i�}�ԊH:R9����"R��T��3��Ԡ#U��ō�Ԡ#U��ŝ���#U��*\D*ϑj Ԍ�"E�q!z�qW������+��W�М��M;L&�EN�k���	}��X�e2!0PK�L&F �i�Ʉ�@c4㲄�@d4㲄�@e4㲄� i!�)+C�q��YA������^�Pb���Z*l�B�BzwJ������ޝS��&*$+�wQT(��
�
o����2�
�u�B�B�_��XHV�8,!/PV�x,�/PVH�L'�
i���@Y!�2��(+�]�e���tBd���qYBe���rj����������|3�7��c�����l.�ݡ_}�����v����� �r��n~h#���=��������vۖk��g�{��LO]��NSm�ol��n������L��h��;��+�ʒ�0!�&�֍EB׌մ�̊c߻�v��u��O�I���{�W��W_���?*[�v�;����Ϯ�]?���M�g��f�����گ�W##,F��92�YTU���n*��9�׏kw16�3i\c�T�4ee-��7�ͩ�vg����1���3ZH��:����
cX��B1m�f��~ �Lg��H����ɑ|~QN]�P�$����ԇGjp����i����kǠ�Fe�����Wem�a��f�]�����*צ�1*DU!�,G�{5�jXm*Ei�S�?�S��
}J���y�ޏ:��C��}�\U�*+�BBY��45ⲩ�W�)ƘkT�V��V�F��q�`T�#�yS[��4�	x���a��ҋZH�8sY�4�W�B6��Ҕ��cQl��2ş}w�������K��BrVplȉ�v��u�|υ,VS�?'c��t��=��}X�u��:m�����wO¥�� �r
�g�^Q]`����;�'�,|�2b�+���>��O/N"ݜR��&�٠�{m��?���6>��J��
 q��\/�oW���������GC��/m��G��є��xt�>e���og��#|2B��F�:�w�F����m���������J�����<Eڳ�h��a!3I�.-=XP��3��f���F�a!s`2��h�{�������� �_TU�_o�����J�E>�~������v�v�߿�����"�MpH�zHké0H5�AJR�LM0���UR%��v�A���l|@ee|A��Ce����/�o������NG`��#D�o(mfS��X��e�aJ��eu��(m�D�g�_?dA���䶬�\�a��%����L#�2����(N?U��@���Ǘ�PK
   � ~X
0�0�  ��                   cirkitFile.jsonPK
   � ~XWC��)�  � /             	  images/093f54e3-331f-4155-80d0-fca9fbcaa25c.pngPK
   JrX�Rr5�  5 /             �  images/1c16f167-bc9c-409e-bb79-de4c62b914f3.pngPK
   � ~X��_8
  3
  /             � images/57489f55-55cc-4ea4-8258-f1cf3d9c722d.pngPK
   � ~X�IM��  � /             �� images/86917e2b-5e70-481a-b4c7-aed39e2d087b.pngPK
   JrX�@M��  2�  /             م images/a3f7833e-13f8-4e96-ad38-aa22696f9742.pngPK
   � ~X`$} [ /             � images/a8bb870d-02b9-45f0-bd60-404fdaa8f6ff.pngPK
   � ~Xp>r�  �  /             J� images/c13bb491-011f-4ad1-adfa-58d33d2d83a5.pngPK
   � ~X�+�s;  z;  /             �� images/f3037bb0-f56a-43e4-a2ff-17056f7c669b.pngPK
   � ~Xϵ��@  �2               O� jsons/user_defined.jsonPK    
 
 j  ��   